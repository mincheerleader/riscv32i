// Verilog netlist created by TD v4.3.815
// Fri Mar 22 14:31:42 2019

`timescale 1ns / 1ps
module __top  // __top.v(3)
  (
  clock,
  rst,
  led
  );

  input clock;  // __top.v(4)
  input rst;  // __top.v(3)
  output led;  // __top.v(5)

  wire [31:0] addr;  // __top.v(17)
  wire [312:0] \cfg_int/wrapper_cfg_inst/reg_inst/cshift_r ;  // D:/td/td/cw\register.v(15)
  wire [17:0] \cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 ;  // D:/td/td/cw\register.v(16)
  wire [31:0] i_data;  // __top.v(15)
  wire [3:0] \m/dram_c0_di ;
  wire [3:0] \m/dram_c0_waddr ;
  wire [3:0] \m/dram_c1_di ;
  wire [3:0] \m/dram_c1_waddr ;
  wire [3:0] \m/dram_c2_di ;
  wire [3:0] \m/dram_c2_waddr ;
  wire [3:0] \m/dram_c3_di ;
  wire [3:0] \m/dram_c3_waddr ;
  wire [3:0] \m/dram_c4_di ;
  wire [3:0] \m/dram_c4_waddr ;
  wire [3:0] \m/dram_c5_di ;
  wire [3:0] \m/dram_c5_waddr ;
  wire [3:0] \m/dram_c6_di ;
  wire [3:0] \m/dram_c6_waddr ;
  wire [3:0] \m/dram_c7_di ;
  wire [3:0] \m/dram_c7_waddr ;
  wire [3:0] n2;
  wire [3:0] n3;
  wire [29:0] n4;
  wire [30:0] n8;
  wire [31:0] o_data;  // __top.v(16)
  wire [31:0] \t/a/EX_A ;  // cpu.v(47)
  wire [31:0] \t/a/EX_B ;  // cpu.v(48)
  wire [2:0] \t/a/EX_fun3 ;  // cpu.v(49)
  wire [6:0] \t/a/EX_fun7 ;  // cpu.v(41)
  wire [31:0] \t/a/EX_memstraddr ;  // cpu.v(38)
  wire [6:0] \t/a/EX_op ;  // cpu.v(42)
  wire [3:0] \t/a/EX_operation ;  // cpu.v(46)
  wire [4:0] \t/a/EX_rd ;  // cpu.v(45)
  wire [31:0] \t/a/EX_regdat1 ;  // cpu.v(39)
  wire [31:0] \t/a/EX_regdat2 ;  // cpu.v(40)
  wire [4:0] \t/a/EX_rs1 ;  // cpu.v(43)
  wire [4:0] \t/a/EX_rs2 ;  // cpu.v(44)
  wire [2:0] \t/a/ID_fun3 ;  // cpu.v(21)
  wire [6:0] \t/a/ID_fun7 ;  // cpu.v(22)
  wire [31:0] \t/a/ID_jump_addr ;  // cpu.v(28)
  wire [31:0] \t/a/ID_jump_regdat1 ;  // cpu.v(29)
  wire [31:0] \t/a/ID_jump_regdat2 ;  // cpu.v(30)
  wire [31:0] \t/a/ID_memstraddr ;  // cpu.v(26)
  wire [6:0] \t/a/ID_op ;  // cpu.v(20)
  wire [4:0] \t/a/ID_rd ;  // cpu.v(23)
  wire [31:0] \t/a/ID_read_dat1 ;  // cpu.v(36)
  wire [31:0] \t/a/ID_read_dat2 ;  // cpu.v(37)
  wire [4:0] \t/a/ID_rs1 ;  // cpu.v(24)
  wire [4:0] \t/a/ID_rs2 ;  // cpu.v(25)
  wire [31:0] \t/a/IF_skip_addr ;  // cpu.v(17)
  wire [31:0] \t/a/MEM_aludat ;  // cpu.v(54)
  wire [2:0] \t/a/MEM_fun3 ;  // cpu.v(58)
  wire [6:0] \t/a/MEM_op ;  // cpu.v(55)
  wire [4:0] \t/a/MEM_rd ;  // cpu.v(56)
  wire [31:0] \t/a/MEM_regdat2 ;  // cpu.v(57)
  wire [6:0] \t/a/WB_op ;  // cpu.v(71)
  wire [4:0] \t/a/WB_rd ;  // cpu.v(70)
  wire  \t/a/alu/mux0_b1/B1_0 ;
  wire  \t/a/alu/mux0_b2/B1_0 ;
  wire  \t/a/alu/mux0_b3/B1_0 ;
  wire  \t/a/alu/mux0_b5/B1_0 ;
  wire  \t/a/alu/mux0_b6/B1_0 ;
  wire [31:0] \t/a/alu/n5 ;
  wire [31:0] \t/a/alu/n6 ;
  wire [1:0] \t/a/alu_A_select ;  // cpu.v(33)
  wire [1:0] \t/a/alu_B_select ;  // cpu.v(34)
  wire [31:0] \t/a/aludat ;  // cpu.v(52)
  wire  \t/a/aluin/sel0_b0/B0 ;
  wire  \t/a/aluin/sel0_b1/B0 ;
  wire  \t/a/aluin/sel0_b10/B0 ;
  wire  \t/a/aluin/sel0_b11/B0 ;
  wire  \t/a/aluin/sel0_b12/B0 ;
  wire  \t/a/aluin/sel0_b13/B0 ;
  wire  \t/a/aluin/sel0_b14/B0 ;
  wire  \t/a/aluin/sel0_b15/B0 ;
  wire  \t/a/aluin/sel0_b16/B0 ;
  wire  \t/a/aluin/sel0_b17/B0 ;
  wire  \t/a/aluin/sel0_b18/B0 ;
  wire  \t/a/aluin/sel0_b19/B0 ;
  wire  \t/a/aluin/sel0_b2/B0 ;
  wire  \t/a/aluin/sel0_b20/B0 ;
  wire  \t/a/aluin/sel0_b21/B0 ;
  wire  \t/a/aluin/sel0_b22/B0 ;
  wire  \t/a/aluin/sel0_b23/B0 ;
  wire  \t/a/aluin/sel0_b24/B0 ;
  wire  \t/a/aluin/sel0_b25/B0 ;
  wire  \t/a/aluin/sel0_b26/B0 ;
  wire  \t/a/aluin/sel0_b27/B0 ;
  wire  \t/a/aluin/sel0_b28/B0 ;
  wire  \t/a/aluin/sel0_b29/B0 ;
  wire  \t/a/aluin/sel0_b3/B0 ;
  wire  \t/a/aluin/sel0_b30/B0 ;
  wire  \t/a/aluin/sel0_b31/B0 ;
  wire  \t/a/aluin/sel0_b4/B0 ;
  wire  \t/a/aluin/sel0_b5/B0 ;
  wire  \t/a/aluin/sel0_b6/B0 ;
  wire  \t/a/aluin/sel0_b7/B0 ;
  wire  \t/a/aluin/sel0_b8/B0 ;
  wire  \t/a/aluin/sel0_b9/B0 ;
  wire  \t/a/aluin/sel1_b10/B9 ;
  wire  \t/a/aluin/sel1_b11/B9 ;
  wire  \t/a/aluin/sel1_b12/B9 ;
  wire  \t/a/aluin/sel1_b13/B9 ;
  wire  \t/a/aluin/sel1_b14/B9 ;
  wire  \t/a/aluin/sel1_b15/B9 ;
  wire  \t/a/aluin/sel1_b16/B9 ;
  wire  \t/a/aluin/sel1_b17/B9 ;
  wire  \t/a/aluin/sel1_b18/B9 ;
  wire  \t/a/aluin/sel1_b19/B9 ;
  wire  \t/a/aluin/sel1_b20/B9 ;
  wire  \t/a/aluin/sel1_b21/B9 ;
  wire  \t/a/aluin/sel1_b22/B9 ;
  wire  \t/a/aluin/sel1_b23/B9 ;
  wire  \t/a/aluin/sel1_b24/B9 ;
  wire  \t/a/aluin/sel1_b25/B9 ;
  wire  \t/a/aluin/sel1_b26/B9 ;
  wire  \t/a/aluin/sel1_b27/B9 ;
  wire  \t/a/aluin/sel1_b28/B9 ;
  wire  \t/a/aluin/sel1_b29/B9 ;
  wire  \t/a/aluin/sel1_b30/B9 ;
  wire  \t/a/aluin/sel1_b31/B9 ;
  wire  \t/a/aluin/sel1_b5/B9 ;
  wire  \t/a/aluin/sel1_b6/B9 ;
  wire  \t/a/aluin/sel1_b7/B9 ;
  wire  \t/a/aluin/sel1_b8/B9 ;
  wire  \t/a/aluin/sel1_b9/B9 ;
  wire [31:0] \t/a/condition/n3 ;
  wire [31:0] \t/a/condition/n5 ;
  wire  \t/a/condition/sel0_b12/B1 ;
  wire  \t/a/condition/sel1/B2 ;
  wire [31:0] \t/a/instr/n12 ;
  wire [29:0] \t/a/instr/n16 ;
  wire  \t/a/mux4_b7/B0_0 ;
  wire [31:0] \t/a/reg_writedat ;  // cpu.v(68)
  wire [31:0] \t/a/regfile/n46 ;
  wire [31:0] \t/a/regfile/regfile$0$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$1$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$10$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$11$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$12$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$13$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$14$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$15$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$16$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$17$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$18$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$19$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$2$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$20$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$21$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$22$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$23$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$24$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$25$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$26$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$27$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$28$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$29$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$3$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$30$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$31$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$4$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$5$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$6$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$7$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$8$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$9$ ;  // register.v(5)
  wire [31:0] \t/busarbitration/instruction ;  // io.v(35)
  wire [31:0] \t/memstraddress ;  // top2.v(17)
  wire [15:0] \trig_node/trigger_node_int_0/force_acq_len ;  // D:/td/td/cw\trigger_node.v(37)
  wire [15:0] \trig_node/trigger_node_int_0/force_acq_reg ;  // D:/td/td/cw\trigger_node.v(39)
  wire [15:0] \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp ;  // D:/td/td/cw\write_ctrl.v(15)
  wire [19:0] \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 ;
  wire [15:0] \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 ;
  wire [15:0] \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 ;
  wire [15:0] \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count ;  // D:/td/td/cw\write_ctrl.v(19)
  wire [16:0] \trig_node/trigger_node_int_0/n141 ;
  wire [15:0] \trig_node/trigger_node_int_0/n179 ;
  wire _al_u1000_o;
  wire _al_u1001_o;
  wire _al_u1002_o;
  wire _al_u1003_o;
  wire _al_u1004_o;
  wire _al_u1043_o;
  wire _al_u1044_o;
  wire _al_u1045_o;
  wire _al_u1046_o;
  wire _al_u1047_o;
  wire _al_u1049_o;
  wire _al_u1050_o;
  wire _al_u1051_o;
  wire _al_u1052_o;
  wire _al_u1053_o;
  wire _al_u1054_o;
  wire _al_u1055_o;
  wire _al_u1056_o;
  wire _al_u1057_o;
  wire _al_u1058_o;
  wire _al_u1059_o;
  wire _al_u1060_o;
  wire _al_u1061_o;
  wire _al_u1062_o;
  wire _al_u1063_o;
  wire _al_u1064_o;
  wire _al_u1065_o;
  wire _al_u1066_o;
  wire _al_u1067_o;
  wire _al_u1068_o;
  wire _al_u1069_o;
  wire _al_u1071_o;
  wire _al_u1072_o;
  wire _al_u1073_o;
  wire _al_u1074_o;
  wire _al_u1075_o;
  wire _al_u1076_o;
  wire _al_u1077_o;
  wire _al_u1078_o;
  wire _al_u1079_o;
  wire _al_u1080_o;
  wire _al_u1081_o;
  wire _al_u1082_o;
  wire _al_u1083_o;
  wire _al_u1084_o;
  wire _al_u1085_o;
  wire _al_u1086_o;
  wire _al_u1087_o;
  wire _al_u1088_o;
  wire _al_u1089_o;
  wire _al_u1090_o;
  wire _al_u1092_o;
  wire _al_u1093_o;
  wire _al_u1094_o;
  wire _al_u1095_o;
  wire _al_u1096_o;
  wire _al_u1097_o;
  wire _al_u1098_o;
  wire _al_u1099_o;
  wire _al_u1100_o;
  wire _al_u1101_o;
  wire _al_u1102_o;
  wire _al_u1103_o;
  wire _al_u1104_o;
  wire _al_u1105_o;
  wire _al_u1106_o;
  wire _al_u1107_o;
  wire _al_u1108_o;
  wire _al_u1109_o;
  wire _al_u1110_o;
  wire _al_u1111_o;
  wire _al_u1113_o;
  wire _al_u1114_o;
  wire _al_u1115_o;
  wire _al_u1116_o;
  wire _al_u1117_o;
  wire _al_u1118_o;
  wire _al_u1119_o;
  wire _al_u1120_o;
  wire _al_u1121_o;
  wire _al_u1122_o;
  wire _al_u1123_o;
  wire _al_u1124_o;
  wire _al_u1125_o;
  wire _al_u1126_o;
  wire _al_u1127_o;
  wire _al_u1128_o;
  wire _al_u1129_o;
  wire _al_u1130_o;
  wire _al_u1131_o;
  wire _al_u1132_o;
  wire _al_u1134_o;
  wire _al_u1135_o;
  wire _al_u1136_o;
  wire _al_u1137_o;
  wire _al_u1138_o;
  wire _al_u1139_o;
  wire _al_u1140_o;
  wire _al_u1141_o;
  wire _al_u1142_o;
  wire _al_u1143_o;
  wire _al_u1144_o;
  wire _al_u1145_o;
  wire _al_u1146_o;
  wire _al_u1147_o;
  wire _al_u1148_o;
  wire _al_u1149_o;
  wire _al_u1150_o;
  wire _al_u1151_o;
  wire _al_u1152_o;
  wire _al_u1153_o;
  wire _al_u1155_o;
  wire _al_u1156_o;
  wire _al_u1157_o;
  wire _al_u1158_o;
  wire _al_u1159_o;
  wire _al_u1160_o;
  wire _al_u1161_o;
  wire _al_u1162_o;
  wire _al_u1163_o;
  wire _al_u1164_o;
  wire _al_u1165_o;
  wire _al_u1166_o;
  wire _al_u1167_o;
  wire _al_u1168_o;
  wire _al_u1169_o;
  wire _al_u1170_o;
  wire _al_u1171_o;
  wire _al_u1172_o;
  wire _al_u1173_o;
  wire _al_u1174_o;
  wire _al_u1176_o;
  wire _al_u1177_o;
  wire _al_u1178_o;
  wire _al_u1179_o;
  wire _al_u1180_o;
  wire _al_u1181_o;
  wire _al_u1182_o;
  wire _al_u1183_o;
  wire _al_u1184_o;
  wire _al_u1185_o;
  wire _al_u1186_o;
  wire _al_u1187_o;
  wire _al_u1188_o;
  wire _al_u1189_o;
  wire _al_u1190_o;
  wire _al_u1191_o;
  wire _al_u1192_o;
  wire _al_u1193_o;
  wire _al_u1194_o;
  wire _al_u1195_o;
  wire _al_u1197_o;
  wire _al_u1198_o;
  wire _al_u1199_o;
  wire _al_u1200_o;
  wire _al_u1201_o;
  wire _al_u1202_o;
  wire _al_u1203_o;
  wire _al_u1204_o;
  wire _al_u1205_o;
  wire _al_u1206_o;
  wire _al_u1207_o;
  wire _al_u1208_o;
  wire _al_u1209_o;
  wire _al_u1210_o;
  wire _al_u1211_o;
  wire _al_u1212_o;
  wire _al_u1213_o;
  wire _al_u1214_o;
  wire _al_u1215_o;
  wire _al_u1216_o;
  wire _al_u1218_o;
  wire _al_u1219_o;
  wire _al_u1220_o;
  wire _al_u1221_o;
  wire _al_u1222_o;
  wire _al_u1223_o;
  wire _al_u1224_o;
  wire _al_u1225_o;
  wire _al_u1226_o;
  wire _al_u1227_o;
  wire _al_u1228_o;
  wire _al_u1229_o;
  wire _al_u1230_o;
  wire _al_u1231_o;
  wire _al_u1232_o;
  wire _al_u1233_o;
  wire _al_u1234_o;
  wire _al_u1235_o;
  wire _al_u1236_o;
  wire _al_u1237_o;
  wire _al_u1239_o;
  wire _al_u1240_o;
  wire _al_u1241_o;
  wire _al_u1242_o;
  wire _al_u1243_o;
  wire _al_u1244_o;
  wire _al_u1245_o;
  wire _al_u1246_o;
  wire _al_u1247_o;
  wire _al_u1248_o;
  wire _al_u1249_o;
  wire _al_u1250_o;
  wire _al_u1251_o;
  wire _al_u1252_o;
  wire _al_u1253_o;
  wire _al_u1254_o;
  wire _al_u1255_o;
  wire _al_u1256_o;
  wire _al_u1257_o;
  wire _al_u1258_o;
  wire _al_u1260_o;
  wire _al_u1261_o;
  wire _al_u1262_o;
  wire _al_u1263_o;
  wire _al_u1264_o;
  wire _al_u1265_o;
  wire _al_u1266_o;
  wire _al_u1267_o;
  wire _al_u1268_o;
  wire _al_u1269_o;
  wire _al_u1270_o;
  wire _al_u1271_o;
  wire _al_u1272_o;
  wire _al_u1273_o;
  wire _al_u1274_o;
  wire _al_u1275_o;
  wire _al_u1276_o;
  wire _al_u1277_o;
  wire _al_u1278_o;
  wire _al_u1279_o;
  wire _al_u1281_o;
  wire _al_u1282_o;
  wire _al_u1283_o;
  wire _al_u1284_o;
  wire _al_u1285_o;
  wire _al_u1286_o;
  wire _al_u1287_o;
  wire _al_u1288_o;
  wire _al_u1289_o;
  wire _al_u1290_o;
  wire _al_u1291_o;
  wire _al_u1292_o;
  wire _al_u1293_o;
  wire _al_u1294_o;
  wire _al_u1295_o;
  wire _al_u1296_o;
  wire _al_u1297_o;
  wire _al_u1298_o;
  wire _al_u1299_o;
  wire _al_u1300_o;
  wire _al_u1302_o;
  wire _al_u1303_o;
  wire _al_u1304_o;
  wire _al_u1305_o;
  wire _al_u1306_o;
  wire _al_u1307_o;
  wire _al_u1308_o;
  wire _al_u1309_o;
  wire _al_u1310_o;
  wire _al_u1311_o;
  wire _al_u1312_o;
  wire _al_u1313_o;
  wire _al_u1314_o;
  wire _al_u1315_o;
  wire _al_u1316_o;
  wire _al_u1317_o;
  wire _al_u1318_o;
  wire _al_u1319_o;
  wire _al_u1320_o;
  wire _al_u1321_o;
  wire _al_u1323_o;
  wire _al_u1324_o;
  wire _al_u1325_o;
  wire _al_u1326_o;
  wire _al_u1327_o;
  wire _al_u1328_o;
  wire _al_u1329_o;
  wire _al_u1330_o;
  wire _al_u1331_o;
  wire _al_u1332_o;
  wire _al_u1333_o;
  wire _al_u1334_o;
  wire _al_u1335_o;
  wire _al_u1336_o;
  wire _al_u1337_o;
  wire _al_u1338_o;
  wire _al_u1339_o;
  wire _al_u1340_o;
  wire _al_u1341_o;
  wire _al_u1342_o;
  wire _al_u1344_o;
  wire _al_u1345_o;
  wire _al_u1346_o;
  wire _al_u1347_o;
  wire _al_u1348_o;
  wire _al_u1349_o;
  wire _al_u1350_o;
  wire _al_u1351_o;
  wire _al_u1352_o;
  wire _al_u1353_o;
  wire _al_u1354_o;
  wire _al_u1355_o;
  wire _al_u1356_o;
  wire _al_u1357_o;
  wire _al_u1358_o;
  wire _al_u1359_o;
  wire _al_u1360_o;
  wire _al_u1361_o;
  wire _al_u1362_o;
  wire _al_u1363_o;
  wire _al_u1365_o;
  wire _al_u1366_o;
  wire _al_u1367_o;
  wire _al_u1368_o;
  wire _al_u1369_o;
  wire _al_u1370_o;
  wire _al_u1371_o;
  wire _al_u1372_o;
  wire _al_u1373_o;
  wire _al_u1374_o;
  wire _al_u1375_o;
  wire _al_u1376_o;
  wire _al_u1377_o;
  wire _al_u1378_o;
  wire _al_u1379_o;
  wire _al_u1380_o;
  wire _al_u1381_o;
  wire _al_u1382_o;
  wire _al_u1383_o;
  wire _al_u1384_o;
  wire _al_u1386_o;
  wire _al_u1387_o;
  wire _al_u1388_o;
  wire _al_u1389_o;
  wire _al_u1390_o;
  wire _al_u1391_o;
  wire _al_u1392_o;
  wire _al_u1393_o;
  wire _al_u1394_o;
  wire _al_u1395_o;
  wire _al_u1396_o;
  wire _al_u1397_o;
  wire _al_u1398_o;
  wire _al_u1399_o;
  wire _al_u1400_o;
  wire _al_u1401_o;
  wire _al_u1402_o;
  wire _al_u1403_o;
  wire _al_u1404_o;
  wire _al_u1405_o;
  wire _al_u1407_o;
  wire _al_u1408_o;
  wire _al_u1409_o;
  wire _al_u1410_o;
  wire _al_u1411_o;
  wire _al_u1412_o;
  wire _al_u1413_o;
  wire _al_u1414_o;
  wire _al_u1415_o;
  wire _al_u1416_o;
  wire _al_u1417_o;
  wire _al_u1418_o;
  wire _al_u1419_o;
  wire _al_u1420_o;
  wire _al_u1421_o;
  wire _al_u1422_o;
  wire _al_u1423_o;
  wire _al_u1424_o;
  wire _al_u1425_o;
  wire _al_u1426_o;
  wire _al_u1428_o;
  wire _al_u1429_o;
  wire _al_u1430_o;
  wire _al_u1431_o;
  wire _al_u1432_o;
  wire _al_u1433_o;
  wire _al_u1434_o;
  wire _al_u1435_o;
  wire _al_u1436_o;
  wire _al_u1437_o;
  wire _al_u1438_o;
  wire _al_u1439_o;
  wire _al_u1440_o;
  wire _al_u1441_o;
  wire _al_u1442_o;
  wire _al_u1443_o;
  wire _al_u1444_o;
  wire _al_u1445_o;
  wire _al_u1446_o;
  wire _al_u1447_o;
  wire _al_u1449_o;
  wire _al_u1450_o;
  wire _al_u1451_o;
  wire _al_u1452_o;
  wire _al_u1453_o;
  wire _al_u1454_o;
  wire _al_u1455_o;
  wire _al_u1456_o;
  wire _al_u1457_o;
  wire _al_u1458_o;
  wire _al_u1459_o;
  wire _al_u1460_o;
  wire _al_u1461_o;
  wire _al_u1462_o;
  wire _al_u1463_o;
  wire _al_u1464_o;
  wire _al_u1465_o;
  wire _al_u1466_o;
  wire _al_u1467_o;
  wire _al_u1468_o;
  wire _al_u1470_o;
  wire _al_u1471_o;
  wire _al_u1472_o;
  wire _al_u1473_o;
  wire _al_u1474_o;
  wire _al_u1475_o;
  wire _al_u1476_o;
  wire _al_u1477_o;
  wire _al_u1478_o;
  wire _al_u1479_o;
  wire _al_u1480_o;
  wire _al_u1481_o;
  wire _al_u1482_o;
  wire _al_u1483_o;
  wire _al_u1484_o;
  wire _al_u1485_o;
  wire _al_u1486_o;
  wire _al_u1487_o;
  wire _al_u1488_o;
  wire _al_u1489_o;
  wire _al_u1491_o;
  wire _al_u1492_o;
  wire _al_u1493_o;
  wire _al_u1494_o;
  wire _al_u1495_o;
  wire _al_u1496_o;
  wire _al_u1497_o;
  wire _al_u1498_o;
  wire _al_u1499_o;
  wire _al_u1500_o;
  wire _al_u1501_o;
  wire _al_u1502_o;
  wire _al_u1503_o;
  wire _al_u1504_o;
  wire _al_u1505_o;
  wire _al_u1506_o;
  wire _al_u1507_o;
  wire _al_u1508_o;
  wire _al_u1509_o;
  wire _al_u1510_o;
  wire _al_u1512_o;
  wire _al_u1513_o;
  wire _al_u1514_o;
  wire _al_u1515_o;
  wire _al_u1516_o;
  wire _al_u1517_o;
  wire _al_u1518_o;
  wire _al_u1519_o;
  wire _al_u1520_o;
  wire _al_u1521_o;
  wire _al_u1522_o;
  wire _al_u1523_o;
  wire _al_u1524_o;
  wire _al_u1525_o;
  wire _al_u1526_o;
  wire _al_u1527_o;
  wire _al_u1528_o;
  wire _al_u1529_o;
  wire _al_u1530_o;
  wire _al_u1531_o;
  wire _al_u1533_o;
  wire _al_u1534_o;
  wire _al_u1535_o;
  wire _al_u1536_o;
  wire _al_u1537_o;
  wire _al_u1538_o;
  wire _al_u1539_o;
  wire _al_u1540_o;
  wire _al_u1541_o;
  wire _al_u1542_o;
  wire _al_u1543_o;
  wire _al_u1544_o;
  wire _al_u1545_o;
  wire _al_u1546_o;
  wire _al_u1547_o;
  wire _al_u1548_o;
  wire _al_u1549_o;
  wire _al_u1550_o;
  wire _al_u1551_o;
  wire _al_u1552_o;
  wire _al_u1554_o;
  wire _al_u1555_o;
  wire _al_u1556_o;
  wire _al_u1557_o;
  wire _al_u1558_o;
  wire _al_u1559_o;
  wire _al_u1560_o;
  wire _al_u1561_o;
  wire _al_u1562_o;
  wire _al_u1563_o;
  wire _al_u1564_o;
  wire _al_u1565_o;
  wire _al_u1566_o;
  wire _al_u1567_o;
  wire _al_u1568_o;
  wire _al_u1569_o;
  wire _al_u1570_o;
  wire _al_u1571_o;
  wire _al_u1572_o;
  wire _al_u1573_o;
  wire _al_u1575_o;
  wire _al_u1576_o;
  wire _al_u1577_o;
  wire _al_u1578_o;
  wire _al_u1579_o;
  wire _al_u1580_o;
  wire _al_u1581_o;
  wire _al_u1582_o;
  wire _al_u1583_o;
  wire _al_u1584_o;
  wire _al_u1585_o;
  wire _al_u1586_o;
  wire _al_u1587_o;
  wire _al_u1588_o;
  wire _al_u1589_o;
  wire _al_u1590_o;
  wire _al_u1591_o;
  wire _al_u1592_o;
  wire _al_u1593_o;
  wire _al_u1594_o;
  wire _al_u1596_o;
  wire _al_u1597_o;
  wire _al_u1598_o;
  wire _al_u1599_o;
  wire _al_u1600_o;
  wire _al_u1601_o;
  wire _al_u1602_o;
  wire _al_u1603_o;
  wire _al_u1604_o;
  wire _al_u1605_o;
  wire _al_u1606_o;
  wire _al_u1607_o;
  wire _al_u1608_o;
  wire _al_u1609_o;
  wire _al_u1610_o;
  wire _al_u1611_o;
  wire _al_u1612_o;
  wire _al_u1613_o;
  wire _al_u1614_o;
  wire _al_u1615_o;
  wire _al_u1617_o;
  wire _al_u1618_o;
  wire _al_u1619_o;
  wire _al_u1620_o;
  wire _al_u1621_o;
  wire _al_u1622_o;
  wire _al_u1623_o;
  wire _al_u1624_o;
  wire _al_u1625_o;
  wire _al_u1626_o;
  wire _al_u1627_o;
  wire _al_u1628_o;
  wire _al_u1629_o;
  wire _al_u1630_o;
  wire _al_u1631_o;
  wire _al_u1632_o;
  wire _al_u1633_o;
  wire _al_u1634_o;
  wire _al_u1635_o;
  wire _al_u1636_o;
  wire _al_u1638_o;
  wire _al_u1639_o;
  wire _al_u1640_o;
  wire _al_u1641_o;
  wire _al_u1642_o;
  wire _al_u1643_o;
  wire _al_u1644_o;
  wire _al_u1645_o;
  wire _al_u1646_o;
  wire _al_u1647_o;
  wire _al_u1648_o;
  wire _al_u1649_o;
  wire _al_u1650_o;
  wire _al_u1651_o;
  wire _al_u1652_o;
  wire _al_u1653_o;
  wire _al_u1654_o;
  wire _al_u1655_o;
  wire _al_u1656_o;
  wire _al_u1657_o;
  wire _al_u1659_o;
  wire _al_u1660_o;
  wire _al_u1661_o;
  wire _al_u1662_o;
  wire _al_u1663_o;
  wire _al_u1664_o;
  wire _al_u1665_o;
  wire _al_u1666_o;
  wire _al_u1667_o;
  wire _al_u1668_o;
  wire _al_u1669_o;
  wire _al_u1670_o;
  wire _al_u1671_o;
  wire _al_u1672_o;
  wire _al_u1673_o;
  wire _al_u1674_o;
  wire _al_u1675_o;
  wire _al_u1676_o;
  wire _al_u1677_o;
  wire _al_u1678_o;
  wire _al_u1680_o;
  wire _al_u1681_o;
  wire _al_u1682_o;
  wire _al_u1683_o;
  wire _al_u1684_o;
  wire _al_u1685_o;
  wire _al_u1686_o;
  wire _al_u1687_o;
  wire _al_u1688_o;
  wire _al_u1689_o;
  wire _al_u1690_o;
  wire _al_u1691_o;
  wire _al_u1692_o;
  wire _al_u1693_o;
  wire _al_u1694_o;
  wire _al_u1695_o;
  wire _al_u1696_o;
  wire _al_u1697_o;
  wire _al_u1698_o;
  wire _al_u1699_o;
  wire _al_u1701_o;
  wire _al_u1702_o;
  wire _al_u1703_o;
  wire _al_u1704_o;
  wire _al_u1705_o;
  wire _al_u1706_o;
  wire _al_u1707_o;
  wire _al_u1708_o;
  wire _al_u1709_o;
  wire _al_u1710_o;
  wire _al_u1711_o;
  wire _al_u1712_o;
  wire _al_u1713_o;
  wire _al_u1714_o;
  wire _al_u1715_o;
  wire _al_u1716_o;
  wire _al_u1717_o;
  wire _al_u1718_o;
  wire _al_u1719_o;
  wire _al_u1720_o;
  wire _al_u1722_o;
  wire _al_u1723_o;
  wire _al_u1724_o;
  wire _al_u1725_o;
  wire _al_u1727_o;
  wire _al_u1728_o;
  wire _al_u1729_o;
  wire _al_u1730_o;
  wire _al_u1733_o;
  wire _al_u1734_o;
  wire _al_u1735_o;
  wire _al_u1736_o;
  wire _al_u1737_o;
  wire _al_u1739_o;
  wire _al_u1740_o;
  wire _al_u1742_o;
  wire _al_u1743_o;
  wire _al_u1744_o;
  wire _al_u1745_o;
  wire _al_u1747_o;
  wire _al_u1783_o;
  wire _al_u1784_o;
  wire _al_u1785_o;
  wire _al_u1786_o;
  wire _al_u1788_o;
  wire _al_u1789_o;
  wire _al_u1790_o;
  wire _al_u1791_o;
  wire _al_u1792_o;
  wire _al_u1793_o;
  wire _al_u1796_o;
  wire _al_u1797_o;
  wire _al_u1798_o;
  wire _al_u1800_o;
  wire _al_u1801_o;
  wire _al_u1802_o;
  wire _al_u1803_o;
  wire _al_u1806_o;
  wire _al_u1808_o;
  wire _al_u1811_o;
  wire _al_u1814_o;
  wire _al_u1817_o;
  wire _al_u1820_o;
  wire _al_u1823_o;
  wire _al_u1826_o;
  wire _al_u1829_o;
  wire _al_u1832_o;
  wire _al_u1835_o;
  wire _al_u1838_o;
  wire _al_u1841_o;
  wire _al_u1844_o;
  wire _al_u1847_o;
  wire _al_u1850_o;
  wire _al_u1853_o;
  wire _al_u1856_o;
  wire _al_u1859_o;
  wire _al_u1862_o;
  wire _al_u1865_o;
  wire _al_u1868_o;
  wire _al_u1871_o;
  wire _al_u1874_o;
  wire _al_u1877_o;
  wire _al_u1880_o;
  wire _al_u1883_o;
  wire _al_u1886_o;
  wire _al_u1889_o;
  wire _al_u1892_o;
  wire _al_u1895_o;
  wire _al_u1898_o;
  wire _al_u1902_o;
  wire _al_u1903_o;
  wire _al_u1904_o;
  wire _al_u1906_o;
  wire _al_u1908_o;
  wire _al_u1916_o;
  wire _al_u1917_o;
  wire _al_u1918_o;
  wire _al_u1935_o;
  wire _al_u1940_o;
  wire _al_u1944_o;
  wire _al_u1947_o;
  wire _al_u1948_o;
  wire _al_u1950_o;
  wire _al_u1956_o;
  wire _al_u1958_o;
  wire _al_u1960_o;
  wire _al_u1962_o;
  wire _al_u1965_o;
  wire _al_u1967_o;
  wire _al_u1968_o;
  wire _al_u1969_o;
  wire _al_u1970_o;
  wire _al_u1973_o;
  wire _al_u1974_o;
  wire _al_u1975_o;
  wire _al_u1976_o;
  wire _al_u1979_o;
  wire _al_u1983_o;
  wire _al_u1984_o;
  wire _al_u1985_o;
  wire _al_u1987_o;
  wire _al_u1990_o;
  wire _al_u1993_o;
  wire _al_u1996_o;
  wire _al_u1999_o;
  wire _al_u2000_o;
  wire _al_u2002_o;
  wire _al_u2005_o;
  wire _al_u2007_o;
  wire _al_u2009_o;
  wire _al_u2010_o;
  wire _al_u2012_o;
  wire _al_u2015_o;
  wire _al_u2018_o;
  wire _al_u2021_o;
  wire _al_u2024_o;
  wire _al_u2027_o;
  wire _al_u2030_o;
  wire _al_u2033_o;
  wire _al_u2036_o;
  wire _al_u2039_o;
  wire _al_u2042_o;
  wire _al_u2045_o;
  wire _al_u2048_o;
  wire _al_u2051_o;
  wire _al_u2054_o;
  wire _al_u2057_o;
  wire _al_u2060_o;
  wire _al_u2063_o;
  wire _al_u2066_o;
  wire _al_u2069_o;
  wire _al_u2072_o;
  wire _al_u2073_o;
  wire _al_u2075_o;
  wire _al_u2076_o;
  wire _al_u2078_o;
  wire _al_u2080_o;
  wire _al_u2092_o;
  wire _al_u2093_o;
  wire _al_u2095_o;
  wire _al_u2096_o;
  wire _al_u2097_o;
  wire _al_u2098_o;
  wire _al_u2099_o;
  wire _al_u2100_o;
  wire _al_u2101_o;
  wire _al_u2102_o;
  wire _al_u2103_o;
  wire _al_u2104_o;
  wire _al_u2105_o;
  wire _al_u2106_o;
  wire _al_u2107_o;
  wire _al_u2109_o;
  wire _al_u2111_o;
  wire _al_u2113_o;
  wire _al_u2115_o;
  wire _al_u2117_o;
  wire _al_u2119_o;
  wire _al_u2124_o;
  wire _al_u2126_o;
  wire _al_u2128_o;
  wire _al_u2130_o;
  wire _al_u2133_o;
  wire _al_u2136_o;
  wire _al_u2137_o;
  wire _al_u2140_o;
  wire _al_u2143_o;
  wire _al_u2144_o;
  wire _al_u2145_o;
  wire _al_u2146_o;
  wire _al_u2147_o;
  wire _al_u2150_o;
  wire _al_u2153_o;
  wire _al_u2154_o;
  wire _al_u2157_o;
  wire _al_u2159_o;
  wire _al_u2161_o;
  wire _al_u2162_o;
  wire _al_u2163_o;
  wire _al_u2165_o;
  wire _al_u2166_o;
  wire _al_u2168_o;
  wire _al_u2169_o;
  wire _al_u2170_o;
  wire _al_u2172_o;
  wire _al_u2175_o;
  wire _al_u2178_o;
  wire _al_u2179_o;
  wire _al_u2182_o;
  wire _al_u2184_o;
  wire _al_u2185_o;
  wire _al_u2186_o;
  wire _al_u2187_o;
  wire _al_u2188_o;
  wire _al_u2191_o;
  wire _al_u2194_o;
  wire _al_u2195_o;
  wire _al_u2198_o;
  wire _al_u2201_o;
  wire _al_u2202_o;
  wire _al_u2203_o;
  wire _al_u2208_o;
  wire _al_u2209_o;
  wire _al_u2210_o;
  wire _al_u2212_o;
  wire _al_u2213_o;
  wire _al_u2214_o;
  wire _al_u2215_o;
  wire _al_u2216_o;
  wire _al_u2218_o;
  wire _al_u2219_o;
  wire _al_u2220_o;
  wire _al_u2221_o;
  wire _al_u2222_o;
  wire _al_u2223_o;
  wire _al_u2224_o;
  wire _al_u2225_o;
  wire _al_u2226_o;
  wire _al_u2227_o;
  wire _al_u2229_o;
  wire _al_u2232_o;
  wire _al_u2233_o;
  wire _al_u2234_o;
  wire _al_u2236_o;
  wire _al_u2237_o;
  wire _al_u2238_o;
  wire _al_u2239_o;
  wire _al_u2240_o;
  wire _al_u2241_o;
  wire _al_u2242_o;
  wire _al_u2243_o;
  wire _al_u2244_o;
  wire _al_u2245_o;
  wire _al_u2246_o;
  wire _al_u2247_o;
  wire _al_u2248_o;
  wire _al_u2249_o;
  wire _al_u2250_o;
  wire _al_u2252_o;
  wire _al_u2255_o;
  wire _al_u2256_o;
  wire _al_u2257_o;
  wire _al_u2259_o;
  wire _al_u2260_o;
  wire _al_u2262_o;
  wire _al_u2263_o;
  wire _al_u2264_o;
  wire _al_u2265_o;
  wire _al_u2266_o;
  wire _al_u2267_o;
  wire _al_u2269_o;
  wire _al_u2270_o;
  wire _al_u2272_o;
  wire _al_u2273_o;
  wire _al_u2274_o;
  wire _al_u2276_o;
  wire _al_u2277_o;
  wire _al_u2279_o;
  wire _al_u2280_o;
  wire _al_u2281_o;
  wire _al_u2282_o;
  wire _al_u2283_o;
  wire _al_u2284_o;
  wire _al_u2286_o;
  wire _al_u2287_o;
  wire _al_u2289_o;
  wire _al_u2290_o;
  wire _al_u2291_o;
  wire _al_u2293_o;
  wire _al_u2294_o;
  wire _al_u2296_o;
  wire _al_u2297_o;
  wire _al_u2298_o;
  wire _al_u2299_o;
  wire _al_u2300_o;
  wire _al_u2301_o;
  wire _al_u2303_o;
  wire _al_u2304_o;
  wire _al_u2306_o;
  wire _al_u2307_o;
  wire _al_u2308_o;
  wire _al_u2310_o;
  wire _al_u2311_o;
  wire _al_u2312_o;
  wire _al_u2313_o;
  wire _al_u2314_o;
  wire _al_u2315_o;
  wire _al_u2316_o;
  wire _al_u2317_o;
  wire _al_u2319_o;
  wire _al_u2320_o;
  wire _al_u2322_o;
  wire _al_u2323_o;
  wire _al_u2324_o;
  wire _al_u2327_o;
  wire _al_u2328_o;
  wire _al_u2329_o;
  wire _al_u2330_o;
  wire _al_u2332_o;
  wire _al_u2333_o;
  wire _al_u2334_o;
  wire _al_u2335_o;
  wire _al_u2336_o;
  wire _al_u2337_o;
  wire _al_u2340_o;
  wire _al_u2341_o;
  wire _al_u2342_o;
  wire _al_u2343_o;
  wire _al_u2345_o;
  wire _al_u2346_o;
  wire _al_u2347_o;
  wire _al_u2348_o;
  wire _al_u2349_o;
  wire _al_u2350_o;
  wire _al_u2353_o;
  wire _al_u2354_o;
  wire _al_u2355_o;
  wire _al_u2356_o;
  wire _al_u2358_o;
  wire _al_u2359_o;
  wire _al_u2360_o;
  wire _al_u2361_o;
  wire _al_u2362_o;
  wire _al_u2363_o;
  wire _al_u2366_o;
  wire _al_u2367_o;
  wire _al_u2368_o;
  wire _al_u2369_o;
  wire _al_u2371_o;
  wire _al_u2372_o;
  wire _al_u2373_o;
  wire _al_u2374_o;
  wire _al_u2375_o;
  wire _al_u2376_o;
  wire _al_u2378_o;
  wire _al_u2380_o;
  wire _al_u2381_o;
  wire _al_u2383_o;
  wire _al_u2384_o;
  wire _al_u2385_o;
  wire _al_u2386_o;
  wire _al_u2387_o;
  wire _al_u2388_o;
  wire _al_u2390_o;
  wire _al_u2392_o;
  wire _al_u2393_o;
  wire _al_u2395_o;
  wire _al_u2396_o;
  wire _al_u2397_o;
  wire _al_u2398_o;
  wire _al_u2399_o;
  wire _al_u2400_o;
  wire _al_u2403_o;
  wire _al_u2404_o;
  wire _al_u2405_o;
  wire _al_u2406_o;
  wire _al_u2408_o;
  wire _al_u2409_o;
  wire _al_u2410_o;
  wire _al_u2411_o;
  wire _al_u2412_o;
  wire _al_u2413_o;
  wire _al_u2415_o;
  wire _al_u2416_o;
  wire _al_u2417_o;
  wire _al_u2418_o;
  wire _al_u2420_o;
  wire _al_u2421_o;
  wire _al_u2422_o;
  wire _al_u2423_o;
  wire _al_u2424_o;
  wire _al_u2425_o;
  wire _al_u2427_o;
  wire _al_u2429_o;
  wire _al_u2430_o;
  wire _al_u2431_o;
  wire _al_u2432_o;
  wire _al_u2433_o;
  wire _al_u2434_o;
  wire _al_u2435_o;
  wire _al_u2436_o;
  wire _al_u2438_o;
  wire _al_u2439_o;
  wire _al_u2440_o;
  wire _al_u2442_o;
  wire _al_u2443_o;
  wire _al_u2444_o;
  wire _al_u2445_o;
  wire _al_u2446_o;
  wire _al_u2448_o;
  wire _al_u2449_o;
  wire _al_u2450_o;
  wire _al_u2452_o;
  wire _al_u2453_o;
  wire _al_u2454_o;
  wire _al_u2455_o;
  wire _al_u2456_o;
  wire _al_u2458_o;
  wire _al_u2459_o;
  wire _al_u2460_o;
  wire _al_u2462_o;
  wire _al_u2463_o;
  wire _al_u2464_o;
  wire _al_u2465_o;
  wire _al_u2466_o;
  wire _al_u2468_o;
  wire _al_u2469_o;
  wire _al_u2470_o;
  wire _al_u2472_o;
  wire _al_u2473_o;
  wire _al_u2474_o;
  wire _al_u2475_o;
  wire _al_u2476_o;
  wire _al_u2478_o;
  wire _al_u2479_o;
  wire _al_u2480_o;
  wire _al_u2482_o;
  wire _al_u2483_o;
  wire _al_u2484_o;
  wire _al_u2485_o;
  wire _al_u2486_o;
  wire _al_u2488_o;
  wire _al_u2489_o;
  wire _al_u2490_o;
  wire _al_u2492_o;
  wire _al_u2493_o;
  wire _al_u2494_o;
  wire _al_u2495_o;
  wire _al_u2496_o;
  wire _al_u2498_o;
  wire _al_u2499_o;
  wire _al_u2500_o;
  wire _al_u2502_o;
  wire _al_u2503_o;
  wire _al_u2504_o;
  wire _al_u2505_o;
  wire _al_u2506_o;
  wire _al_u2508_o;
  wire _al_u2509_o;
  wire _al_u2510_o;
  wire _al_u2512_o;
  wire _al_u2513_o;
  wire _al_u2514_o;
  wire _al_u2515_o;
  wire _al_u2516_o;
  wire _al_u251_o;
  wire _al_u2520_o;
  wire _al_u2521_o;
  wire _al_u2522_o;
  wire _al_u2523_o;
  wire _al_u2524_o;
  wire _al_u2525_o;
  wire _al_u2526_o;
  wire _al_u252_o;
  wire _al_u2530_o;
  wire _al_u2531_o;
  wire _al_u2532_o;
  wire _al_u2533_o;
  wire _al_u2534_o;
  wire _al_u2535_o;
  wire _al_u2536_o;
  wire _al_u2538_o;
  wire _al_u2539_o;
  wire _al_u2540_o;
  wire _al_u2541_o;
  wire _al_u2543_o;
  wire _al_u2544_o;
  wire _al_u2545_o;
  wire _al_u2546_o;
  wire _al_u2547_o;
  wire _al_u254_o;
  wire _al_u2551_o;
  wire _al_u2552_o;
  wire _al_u2553_o;
  wire _al_u2554_o;
  wire _al_u2555_o;
  wire _al_u2556_o;
  wire _al_u2560_o;
  wire _al_u2561_o;
  wire _al_u2562_o;
  wire _al_u2563_o;
  wire _al_u2564_o;
  wire _al_u2565_o;
  wire _al_u2567_o;
  wire _al_u2568_o;
  wire _al_u2569_o;
  wire _al_u256_o;
  wire _al_u2570_o;
  wire _al_u2571_o;
  wire _al_u2572_o;
  wire _al_u2573_o;
  wire _al_u2574_o;
  wire _al_u2575_o;
  wire _al_u2576_o;
  wire _al_u2577_o;
  wire _al_u2580_o;
  wire _al_u2581_o;
  wire _al_u2582_o;
  wire _al_u2583_o;
  wire _al_u2584_o;
  wire _al_u2585_o;
  wire _al_u2586_o;
  wire _al_u2587_o;
  wire _al_u2589_o;
  wire _al_u2590_o;
  wire _al_u2591_o;
  wire _al_u2592_o;
  wire _al_u2593_o;
  wire _al_u2594_o;
  wire _al_u2595_o;
  wire _al_u2596_o;
  wire _al_u2597_o;
  wire _al_u2598_o;
  wire _al_u2599_o;
  wire _al_u2600_o;
  wire _al_u2601_o;
  wire _al_u2602_o;
  wire _al_u2604_o;
  wire _al_u2606_o;
  wire _al_u2606_o_placeOpt_1;
  wire _al_u2606_o_placeOpt_2;
  wire _al_u2606_o_placeOpt_3;
  wire _al_u2607_o;
  wire _al_u2608_o;
  wire _al_u2609_o;
  wire _al_u2610_o;
  wire _al_u2610_o_placeOpt_1;
  wire _al_u2610_o_placeOpt_2;
  wire _al_u2610_o_placeOpt_3;
  wire _al_u2611_o;
  wire _al_u2613_o;
  wire _al_u2614_o;
  wire _al_u2614_o_placeOpt_1;
  wire _al_u2614_o_placeOpt_2;
  wire _al_u2614_o_placeOpt_3;
  wire _al_u2615_o;
  wire _al_u2616_o;
  wire _al_u2616_o_placeOpt_1;
  wire _al_u2616_o_placeOpt_2;
  wire _al_u2616_o_placeOpt_3;
  wire _al_u2617_o;
  wire _al_u2619_o;
  wire _al_u2621_o;
  wire _al_u2623_o;
  wire _al_u2625_o;
  wire _al_u2627_o;
  wire _al_u2629_o;
  wire _al_u2631_o;
  wire _al_u2633_o;
  wire _al_u2635_o;
  wire _al_u2637_o;
  wire _al_u2639_o;
  wire _al_u2641_o;
  wire _al_u2643_o;
  wire _al_u2645_o;
  wire _al_u2647_o;
  wire _al_u2649_o;
  wire _al_u2651_o;
  wire _al_u2653_o;
  wire _al_u2655_o;
  wire _al_u2657_o;
  wire _al_u2659_o;
  wire _al_u2661_o;
  wire _al_u2663_o;
  wire _al_u2665_o;
  wire _al_u2667_o;
  wire _al_u2669_o;
  wire _al_u2671_o;
  wire _al_u2673_o;
  wire _al_u2675_o;
  wire _al_u2677_o;
  wire _al_u2679_o;
  wire _al_u2680_o;
  wire _al_u2681_o;
  wire _al_u2683_o;
  wire _al_u2684_o;
  wire _al_u2686_o;
  wire _al_u2687_o;
  wire _al_u2688_o;
  wire _al_u2689_o;
  wire _al_u2690_o;
  wire _al_u2692_o;
  wire _al_u2693_o;
  wire _al_u2695_o;
  wire _al_u2697_o;
  wire _al_u2699_o;
  wire _al_u2701_o;
  wire _al_u2703_o;
  wire _al_u2705_o;
  wire _al_u2707_o;
  wire _al_u2708_o;
  wire _al_u2709_o;
  wire _al_u2710_o;
  wire _al_u2711_o;
  wire _al_u2713_o;
  wire _al_u2714_o;
  wire _al_u2716_o;
  wire _al_u2718_o;
  wire _al_u2720_o;
  wire _al_u2722_o;
  wire _al_u2724_o;
  wire _al_u2726_o;
  wire _al_u2728_o;
  wire _al_u2729_o;
  wire _al_u2730_o;
  wire _al_u2732_o;
  wire _al_u2733_o;
  wire _al_u2735_o;
  wire _al_u2736_o;
  wire _al_u2737_o;
  wire _al_u2739_o;
  wire _al_u2740_o;
  wire _al_u2742_o;
  wire _al_u2744_o;
  wire _al_u2745_o;
  wire _al_u2747_o;
  wire _al_u2748_o;
  wire _al_u2749_o;
  wire _al_u2751_o;
  wire _al_u2752_o;
  wire _al_u2754_o;
  wire _al_u2756_o;
  wire _al_u2758_o;
  wire _al_u2760_o;
  wire _al_u2762_o;
  wire _al_u2764_o;
  wire _al_u2766_o;
  wire _al_u2767_o;
  wire _al_u2768_o;
  wire _al_u2769_o;
  wire _al_u2770_o;
  wire _al_u2771_o;
  wire _al_u2772_o;
  wire _al_u2773_o;
  wire _al_u2774_o;
  wire _al_u2775_o;
  wire _al_u2776_o;
  wire _al_u2777_o;
  wire _al_u2778_o;
  wire _al_u2779_o;
  wire _al_u2780_o;
  wire _al_u2781_o;
  wire _al_u2782_o;
  wire _al_u2783_o;
  wire _al_u2784_o;
  wire _al_u2785_o;
  wire _al_u2786_o;
  wire _al_u2787_o;
  wire _al_u2788_o;
  wire _al_u2789_o;
  wire _al_u2790_o;
  wire _al_u2791_o;
  wire _al_u2792_o;
  wire _al_u2793_o;
  wire _al_u2794_o;
  wire _al_u2795_o;
  wire _al_u2796_o;
  wire _al_u2798_o;
  wire _al_u2799_o;
  wire _al_u2800_o;
  wire _al_u2801_o;
  wire _al_u2802_o;
  wire _al_u2803_o;
  wire _al_u2806_o;
  wire _al_u2807_o;
  wire _al_u2808_o;
  wire _al_u2810_o;
  wire _al_u2811_o;
  wire _al_u2812_o;
  wire _al_u2814_o;
  wire _al_u2815_o;
  wire _al_u2817_o;
  wire _al_u2819_o;
  wire _al_u2821_o;
  wire _al_u2822_o;
  wire _al_u2824_o;
  wire _al_u2826_o;
  wire _al_u2828_o;
  wire _al_u2829_o;
  wire _al_u2831_o;
  wire _al_u2833_o;
  wire _al_u2834_o;
  wire _al_u2836_o;
  wire _al_u2838_o;
  wire _al_u2840_o;
  wire _al_u2841_o;
  wire _al_u2843_o;
  wire _al_u2844_o;
  wire _al_u2846_o;
  wire _al_u2847_o;
  wire _al_u2849_o;
  wire _al_u2850_o;
  wire _al_u2852_o;
  wire _al_u2854_o;
  wire _al_u2856_o;
  wire _al_u2857_o;
  wire _al_u2859_o;
  wire _al_u2860_o;
  wire _al_u2862_o;
  wire _al_u2864_o;
  wire _al_u2866_o;
  wire _al_u2868_o;
  wire _al_u2869_o;
  wire _al_u2871_o;
  wire _al_u2872_o;
  wire _al_u2874_o;
  wire _al_u2875_o;
  wire _al_u2877_o;
  wire _al_u2878_o;
  wire _al_u2880_o;
  wire _al_u2882_o;
  wire _al_u2883_o;
  wire _al_u2885_o;
  wire _al_u2887_o;
  wire _al_u2888_o;
  wire _al_u2890_o;
  wire _al_u290_o;
  wire _al_u3034_o;
  wire _al_u3035_o;
  wire _al_u3055_o;
  wire _al_u3056_o;
  wire _al_u3057_o;
  wire _al_u3058_o;
  wire _al_u3059_o;
  wire _al_u3060_o;
  wire _al_u3061_o;
  wire _al_u3062_o;
  wire _al_u3063_o;
  wire _al_u3064_o;
  wire _al_u3065_o;
  wire _al_u3066_o;
  wire _al_u3067_o;
  wire _al_u3068_o;
  wire _al_u3069_o;
  wire _al_u3071_o;
  wire _al_u3072_o;
  wire _al_u3073_o;
  wire _al_u3074_o;
  wire _al_u3075_o;
  wire _al_u3076_o;
  wire _al_u3077_o;
  wire _al_u3078_o;
  wire _al_u3079_o;
  wire _al_u3080_o;
  wire _al_u3081_o;
  wire _al_u3082_o;
  wire _al_u3083_o;
  wire _al_u3084_o;
  wire _al_u3085_o;
  wire _al_u3086_o;
  wire _al_u3104_o;
  wire _al_u3105_o;
  wire _al_u3106_o;
  wire _al_u3107_o;
  wire _al_u3108_o;
  wire _al_u3109_o;
  wire _al_u3110_o;
  wire _al_u3111_o;
  wire _al_u3112_o;
  wire _al_u3113_o;
  wire _al_u3114_o;
  wire _al_u3115_o;
  wire _al_u3116_o;
  wire _al_u3117_o;
  wire _al_u3118_o;
  wire _al_u3119_o;
  wire _al_u3120_o;
  wire _al_u3121_o;
  wire _al_u3122_o;
  wire _al_u3123_o;
  wire _al_u3124_o;
  wire _al_u3125_o;
  wire _al_u3126_o;
  wire _al_u3127_o;
  wire _al_u3128_o;
  wire _al_u3129_o;
  wire _al_u3130_o;
  wire _al_u3131_o;
  wire _al_u3132_o;
  wire _al_u3133_o;
  wire _al_u3134_o;
  wire _al_u3135_o;
  wire _al_u3136_o;
  wire _al_u3137_o;
  wire _al_u3138_o;
  wire _al_u3139_o;
  wire _al_u3140_o;
  wire _al_u3141_o;
  wire _al_u3142_o;
  wire _al_u3143_o;
  wire _al_u3144_o;
  wire _al_u3145_o;
  wire _al_u3146_o;
  wire _al_u3147_o;
  wire _al_u3148_o;
  wire _al_u3149_o;
  wire _al_u3150_o;
  wire _al_u3151_o;
  wire _al_u3152_o;
  wire _al_u3153_o;
  wire _al_u3154_o;
  wire _al_u3155_o;
  wire _al_u3156_o;
  wire _al_u3157_o;
  wire _al_u3158_o;
  wire _al_u3159_o;
  wire _al_u3160_o;
  wire _al_u3161_o;
  wire _al_u3162_o;
  wire _al_u3163_o;
  wire _al_u3164_o;
  wire _al_u3165_o;
  wire _al_u3166_o;
  wire _al_u3167_o;
  wire _al_u3168_o;
  wire _al_u3169_o;
  wire _al_u3170_o;
  wire _al_u3171_o;
  wire _al_u3172_o;
  wire _al_u3173_o;
  wire _al_u3174_o;
  wire _al_u3175_o;
  wire _al_u3176_o;
  wire _al_u3177_o;
  wire _al_u3178_o;
  wire _al_u3179_o;
  wire _al_u3180_o;
  wire _al_u3181_o;
  wire _al_u3182_o;
  wire _al_u3183_o;
  wire _al_u3184_o;
  wire _al_u3185_o;
  wire _al_u3186_o;
  wire _al_u3187_o;
  wire _al_u3188_o;
  wire _al_u3189_o;
  wire _al_u3190_o;
  wire _al_u3191_o;
  wire _al_u3192_o;
  wire _al_u3193_o;
  wire _al_u3194_o;
  wire _al_u3195_o;
  wire _al_u3196_o;
  wire _al_u3197_o;
  wire _al_u3198_o;
  wire _al_u3199_o;
  wire _al_u3200_o;
  wire _al_u3201_o;
  wire _al_u3202_o;
  wire _al_u3203_o;
  wire _al_u3204_o;
  wire _al_u3205_o;
  wire _al_u3206_o;
  wire _al_u3207_o;
  wire _al_u3208_o;
  wire _al_u3209_o;
  wire _al_u3210_o;
  wire _al_u3211_o;
  wire _al_u3212_o;
  wire _al_u3213_o;
  wire _al_u3214_o;
  wire _al_u3215_o;
  wire _al_u3216_o;
  wire _al_u3217_o;
  wire _al_u3218_o;
  wire _al_u3219_o;
  wire _al_u3220_o;
  wire _al_u3221_o;
  wire _al_u3222_o;
  wire _al_u3223_o;
  wire _al_u3224_o;
  wire _al_u3225_o;
  wire _al_u3226_o;
  wire _al_u3227_o;
  wire _al_u3228_o;
  wire _al_u3229_o;
  wire _al_u3230_o;
  wire _al_u3231_o;
  wire _al_u3232_o;
  wire _al_u3233_o;
  wire _al_u3234_o;
  wire _al_u3235_o;
  wire _al_u3236_o;
  wire _al_u3237_o;
  wire _al_u3238_o;
  wire _al_u3239_o;
  wire _al_u3240_o;
  wire _al_u3241_o;
  wire _al_u3242_o;
  wire _al_u3243_o;
  wire _al_u3244_o;
  wire _al_u3245_o;
  wire _al_u3246_o;
  wire _al_u3247_o;
  wire _al_u3248_o;
  wire _al_u3249_o;
  wire _al_u3250_o;
  wire _al_u3251_o;
  wire _al_u3252_o;
  wire _al_u3253_o;
  wire _al_u3254_o;
  wire _al_u3255_o;
  wire _al_u3256_o;
  wire _al_u3257_o;
  wire _al_u3258_o;
  wire _al_u3259_o;
  wire _al_u3260_o;
  wire _al_u3261_o;
  wire _al_u3262_o;
  wire _al_u3263_o;
  wire _al_u3264_o;
  wire _al_u3265_o;
  wire _al_u3266_o;
  wire _al_u3267_o;
  wire _al_u3268_o;
  wire _al_u3269_o;
  wire _al_u3270_o;
  wire _al_u3271_o;
  wire _al_u3272_o;
  wire _al_u3273_o;
  wire _al_u3274_o;
  wire _al_u3275_o;
  wire _al_u3276_o;
  wire _al_u3277_o;
  wire _al_u3278_o;
  wire _al_u3279_o;
  wire _al_u3280_o;
  wire _al_u3281_o;
  wire _al_u3282_o;
  wire _al_u3283_o;
  wire _al_u3284_o;
  wire _al_u3285_o;
  wire _al_u3286_o;
  wire _al_u3287_o;
  wire _al_u3288_o;
  wire _al_u3289_o;
  wire _al_u328_o;
  wire _al_u3290_o;
  wire _al_u3291_o;
  wire _al_u3292_o;
  wire _al_u3293_o;
  wire _al_u3294_o;
  wire _al_u3295_o;
  wire _al_u3296_o;
  wire _al_u3297_o;
  wire _al_u3298_o;
  wire _al_u3299_o;
  wire _al_u329_o;
  wire _al_u3300_o;
  wire _al_u3301_o;
  wire _al_u3302_o;
  wire _al_u3303_o;
  wire _al_u3304_o;
  wire _al_u3305_o;
  wire _al_u3306_o;
  wire _al_u3307_o;
  wire _al_u3308_o;
  wire _al_u3309_o;
  wire _al_u330_o;
  wire _al_u3310_o;
  wire _al_u3311_o;
  wire _al_u3312_o;
  wire _al_u3313_o;
  wire _al_u3314_o;
  wire _al_u3315_o;
  wire _al_u3316_o;
  wire _al_u3317_o;
  wire _al_u3318_o;
  wire _al_u3319_o;
  wire _al_u331_o;
  wire _al_u3320_o;
  wire _al_u3321_o;
  wire _al_u3322_o;
  wire _al_u3323_o;
  wire _al_u3324_o;
  wire _al_u3325_o;
  wire _al_u3326_o;
  wire _al_u3327_o;
  wire _al_u3328_o;
  wire _al_u3329_o;
  wire _al_u3330_o;
  wire _al_u3331_o;
  wire _al_u3332_o;
  wire _al_u3333_o;
  wire _al_u3334_o;
  wire _al_u3335_o;
  wire _al_u3336_o;
  wire _al_u3337_o;
  wire _al_u3338_o;
  wire _al_u3339_o;
  wire _al_u333_o;
  wire _al_u3340_o;
  wire _al_u3341_o;
  wire _al_u3342_o;
  wire _al_u3343_o;
  wire _al_u3344_o;
  wire _al_u3345_o;
  wire _al_u3346_o;
  wire _al_u3347_o;
  wire _al_u3348_o;
  wire _al_u3349_o;
  wire _al_u334_o;
  wire _al_u3350_o;
  wire _al_u3351_o;
  wire _al_u3352_o;
  wire _al_u3353_o;
  wire _al_u3354_o;
  wire _al_u3355_o;
  wire _al_u3356_o;
  wire _al_u3357_o;
  wire _al_u3358_o;
  wire _al_u3359_o;
  wire _al_u335_o;
  wire _al_u3360_o;
  wire _al_u3361_o;
  wire _al_u3362_o;
  wire _al_u3363_o;
  wire _al_u3364_o;
  wire _al_u3365_o;
  wire _al_u3366_o;
  wire _al_u3367_o;
  wire _al_u3368_o;
  wire _al_u3369_o;
  wire _al_u336_o;
  wire _al_u3370_o;
  wire _al_u3371_o;
  wire _al_u3372_o;
  wire _al_u3373_o;
  wire _al_u3374_o;
  wire _al_u3375_o;
  wire _al_u3376_o;
  wire _al_u3377_o;
  wire _al_u3378_o;
  wire _al_u3379_o;
  wire _al_u337_o;
  wire _al_u3380_o;
  wire _al_u3381_o;
  wire _al_u3382_o;
  wire _al_u3383_o;
  wire _al_u3384_o;
  wire _al_u3385_o;
  wire _al_u3386_o;
  wire _al_u3387_o;
  wire _al_u3388_o;
  wire _al_u3389_o;
  wire _al_u338_o;
  wire _al_u3390_o;
  wire _al_u3391_o;
  wire _al_u3392_o;
  wire _al_u3393_o;
  wire _al_u3394_o;
  wire _al_u3395_o;
  wire _al_u3396_o;
  wire _al_u3397_o;
  wire _al_u3398_o;
  wire _al_u3399_o;
  wire _al_u339_o;
  wire _al_u3400_o;
  wire _al_u3401_o;
  wire _al_u3402_o;
  wire _al_u3403_o;
  wire _al_u3404_o;
  wire _al_u3405_o;
  wire _al_u3406_o;
  wire _al_u3407_o;
  wire _al_u3408_o;
  wire _al_u3409_o;
  wire _al_u340_o;
  wire _al_u3410_o;
  wire _al_u3411_o;
  wire _al_u3412_o;
  wire _al_u3413_o;
  wire _al_u3414_o;
  wire _al_u3415_o;
  wire _al_u3416_o;
  wire _al_u3417_o;
  wire _al_u3418_o;
  wire _al_u3419_o;
  wire _al_u341_o;
  wire _al_u3420_o;
  wire _al_u3421_o;
  wire _al_u3422_o;
  wire _al_u3423_o;
  wire _al_u3424_o;
  wire _al_u3425_o;
  wire _al_u3426_o;
  wire _al_u3427_o;
  wire _al_u3428_o;
  wire _al_u3429_o;
  wire _al_u342_o;
  wire _al_u3430_o;
  wire _al_u3431_o;
  wire _al_u3432_o;
  wire _al_u3433_o;
  wire _al_u3434_o;
  wire _al_u3435_o;
  wire _al_u3436_o;
  wire _al_u3437_o;
  wire _al_u3438_o;
  wire _al_u3439_o;
  wire _al_u343_o;
  wire _al_u3440_o;
  wire _al_u3441_o;
  wire _al_u3442_o;
  wire _al_u3443_o;
  wire _al_u3444_o;
  wire _al_u3445_o;
  wire _al_u3446_o;
  wire _al_u3447_o;
  wire _al_u3448_o;
  wire _al_u3449_o;
  wire _al_u344_o;
  wire _al_u3450_o;
  wire _al_u3451_o;
  wire _al_u3452_o;
  wire _al_u3453_o;
  wire _al_u3454_o;
  wire _al_u3455_o;
  wire _al_u3456_o;
  wire _al_u3457_o;
  wire _al_u3458_o;
  wire _al_u3459_o;
  wire _al_u345_o;
  wire _al_u3460_o;
  wire _al_u3461_o;
  wire _al_u3462_o;
  wire _al_u3463_o;
  wire _al_u3464_o;
  wire _al_u3465_o;
  wire _al_u3466_o;
  wire _al_u3467_o;
  wire _al_u3468_o;
  wire _al_u3469_o;
  wire _al_u346_o;
  wire _al_u3470_o;
  wire _al_u3471_o;
  wire _al_u3472_o;
  wire _al_u3473_o;
  wire _al_u3474_o;
  wire _al_u3475_o;
  wire _al_u3476_o;
  wire _al_u3477_o;
  wire _al_u3478_o;
  wire _al_u3479_o;
  wire _al_u347_o;
  wire _al_u3480_o;
  wire _al_u3481_o;
  wire _al_u3482_o;
  wire _al_u3483_o;
  wire _al_u3484_o;
  wire _al_u3485_o;
  wire _al_u3486_o;
  wire _al_u3487_o;
  wire _al_u3488_o;
  wire _al_u3489_o;
  wire _al_u348_o;
  wire _al_u3490_o;
  wire _al_u3491_o;
  wire _al_u3492_o;
  wire _al_u3493_o;
  wire _al_u3494_o;
  wire _al_u3495_o;
  wire _al_u3496_o;
  wire _al_u3497_o;
  wire _al_u3498_o;
  wire _al_u3499_o;
  wire _al_u349_o;
  wire _al_u3500_o;
  wire _al_u3501_o;
  wire _al_u3502_o;
  wire _al_u3503_o;
  wire _al_u3504_o;
  wire _al_u3505_o;
  wire _al_u3506_o;
  wire _al_u3507_o;
  wire _al_u3508_o;
  wire _al_u3509_o;
  wire _al_u350_o;
  wire _al_u3510_o;
  wire _al_u3511_o;
  wire _al_u3512_o;
  wire _al_u3513_o;
  wire _al_u3514_o;
  wire _al_u3515_o;
  wire _al_u3516_o;
  wire _al_u3517_o;
  wire _al_u3518_o;
  wire _al_u3519_o;
  wire _al_u351_o;
  wire _al_u3520_o;
  wire _al_u3521_o;
  wire _al_u3522_o;
  wire _al_u3523_o;
  wire _al_u3524_o;
  wire _al_u3525_o;
  wire _al_u3526_o;
  wire _al_u3527_o;
  wire _al_u3528_o;
  wire _al_u3529_o;
  wire _al_u352_o;
  wire _al_u3530_o;
  wire _al_u3531_o;
  wire _al_u3532_o;
  wire _al_u3533_o;
  wire _al_u3534_o;
  wire _al_u3535_o;
  wire _al_u3536_o;
  wire _al_u3537_o;
  wire _al_u3538_o;
  wire _al_u3539_o;
  wire _al_u353_o;
  wire _al_u3540_o;
  wire _al_u3541_o;
  wire _al_u3542_o;
  wire _al_u3543_o;
  wire _al_u3544_o;
  wire _al_u3545_o;
  wire _al_u3546_o;
  wire _al_u3547_o;
  wire _al_u355_o;
  wire _al_u356_o;
  wire _al_u357_o;
  wire _al_u358_o;
  wire _al_u359_o;
  wire _al_u360_o;
  wire _al_u361_o;
  wire _al_u362_o;
  wire _al_u363_o;
  wire _al_u364_o;
  wire _al_u365_o;
  wire _al_u366_o;
  wire _al_u367_o;
  wire _al_u368_o;
  wire _al_u369_o;
  wire _al_u370_o;
  wire _al_u371_o;
  wire _al_u372_o;
  wire _al_u373_o;
  wire _al_u374_o;
  wire _al_u376_o;
  wire _al_u377_o;
  wire _al_u378_o;
  wire _al_u379_o;
  wire _al_u380_o;
  wire _al_u381_o;
  wire _al_u382_o;
  wire _al_u383_o;
  wire _al_u384_o;
  wire _al_u385_o;
  wire _al_u386_o;
  wire _al_u387_o;
  wire _al_u388_o;
  wire _al_u389_o;
  wire _al_u390_o;
  wire _al_u391_o;
  wire _al_u392_o;
  wire _al_u393_o;
  wire _al_u394_o;
  wire _al_u395_o;
  wire _al_u397_o;
  wire _al_u398_o;
  wire _al_u399_o;
  wire _al_u400_o;
  wire _al_u401_o;
  wire _al_u402_o;
  wire _al_u403_o;
  wire _al_u404_o;
  wire _al_u405_o;
  wire _al_u406_o;
  wire _al_u407_o;
  wire _al_u408_o;
  wire _al_u409_o;
  wire _al_u410_o;
  wire _al_u411_o;
  wire _al_u412_o;
  wire _al_u413_o;
  wire _al_u414_o;
  wire _al_u415_o;
  wire _al_u416_o;
  wire _al_u418_o;
  wire _al_u419_o;
  wire _al_u420_o;
  wire _al_u421_o;
  wire _al_u422_o;
  wire _al_u423_o;
  wire _al_u424_o;
  wire _al_u425_o;
  wire _al_u426_o;
  wire _al_u427_o;
  wire _al_u428_o;
  wire _al_u429_o;
  wire _al_u430_o;
  wire _al_u431_o;
  wire _al_u432_o;
  wire _al_u433_o;
  wire _al_u434_o;
  wire _al_u435_o;
  wire _al_u436_o;
  wire _al_u437_o;
  wire _al_u439_o;
  wire _al_u440_o;
  wire _al_u441_o;
  wire _al_u442_o;
  wire _al_u443_o;
  wire _al_u444_o;
  wire _al_u445_o;
  wire _al_u446_o;
  wire _al_u447_o;
  wire _al_u448_o;
  wire _al_u449_o;
  wire _al_u450_o;
  wire _al_u451_o;
  wire _al_u452_o;
  wire _al_u453_o;
  wire _al_u454_o;
  wire _al_u455_o;
  wire _al_u456_o;
  wire _al_u457_o;
  wire _al_u458_o;
  wire _al_u460_o;
  wire _al_u461_o;
  wire _al_u462_o;
  wire _al_u463_o;
  wire _al_u464_o;
  wire _al_u465_o;
  wire _al_u466_o;
  wire _al_u467_o;
  wire _al_u468_o;
  wire _al_u469_o;
  wire _al_u470_o;
  wire _al_u471_o;
  wire _al_u472_o;
  wire _al_u473_o;
  wire _al_u474_o;
  wire _al_u475_o;
  wire _al_u476_o;
  wire _al_u477_o;
  wire _al_u478_o;
  wire _al_u479_o;
  wire _al_u481_o;
  wire _al_u482_o;
  wire _al_u483_o;
  wire _al_u484_o;
  wire _al_u485_o;
  wire _al_u486_o;
  wire _al_u487_o;
  wire _al_u488_o;
  wire _al_u489_o;
  wire _al_u490_o;
  wire _al_u491_o;
  wire _al_u492_o;
  wire _al_u493_o;
  wire _al_u494_o;
  wire _al_u495_o;
  wire _al_u496_o;
  wire _al_u497_o;
  wire _al_u498_o;
  wire _al_u499_o;
  wire _al_u500_o;
  wire _al_u502_o;
  wire _al_u503_o;
  wire _al_u504_o;
  wire _al_u505_o;
  wire _al_u506_o;
  wire _al_u507_o;
  wire _al_u508_o;
  wire _al_u509_o;
  wire _al_u510_o;
  wire _al_u511_o;
  wire _al_u512_o;
  wire _al_u513_o;
  wire _al_u514_o;
  wire _al_u515_o;
  wire _al_u516_o;
  wire _al_u517_o;
  wire _al_u518_o;
  wire _al_u519_o;
  wire _al_u520_o;
  wire _al_u521_o;
  wire _al_u523_o;
  wire _al_u524_o;
  wire _al_u525_o;
  wire _al_u526_o;
  wire _al_u527_o;
  wire _al_u528_o;
  wire _al_u529_o;
  wire _al_u530_o;
  wire _al_u531_o;
  wire _al_u532_o;
  wire _al_u533_o;
  wire _al_u534_o;
  wire _al_u535_o;
  wire _al_u536_o;
  wire _al_u537_o;
  wire _al_u538_o;
  wire _al_u539_o;
  wire _al_u540_o;
  wire _al_u541_o;
  wire _al_u542_o;
  wire _al_u544_o;
  wire _al_u545_o;
  wire _al_u546_o;
  wire _al_u547_o;
  wire _al_u548_o;
  wire _al_u549_o;
  wire _al_u550_o;
  wire _al_u551_o;
  wire _al_u552_o;
  wire _al_u553_o;
  wire _al_u554_o;
  wire _al_u555_o;
  wire _al_u556_o;
  wire _al_u557_o;
  wire _al_u558_o;
  wire _al_u559_o;
  wire _al_u560_o;
  wire _al_u561_o;
  wire _al_u562_o;
  wire _al_u563_o;
  wire _al_u565_o;
  wire _al_u566_o;
  wire _al_u567_o;
  wire _al_u568_o;
  wire _al_u569_o;
  wire _al_u570_o;
  wire _al_u571_o;
  wire _al_u572_o;
  wire _al_u573_o;
  wire _al_u574_o;
  wire _al_u575_o;
  wire _al_u576_o;
  wire _al_u577_o;
  wire _al_u578_o;
  wire _al_u579_o;
  wire _al_u580_o;
  wire _al_u581_o;
  wire _al_u582_o;
  wire _al_u583_o;
  wire _al_u584_o;
  wire _al_u586_o;
  wire _al_u587_o;
  wire _al_u588_o;
  wire _al_u589_o;
  wire _al_u590_o;
  wire _al_u591_o;
  wire _al_u592_o;
  wire _al_u593_o;
  wire _al_u594_o;
  wire _al_u595_o;
  wire _al_u596_o;
  wire _al_u597_o;
  wire _al_u598_o;
  wire _al_u599_o;
  wire _al_u600_o;
  wire _al_u601_o;
  wire _al_u602_o;
  wire _al_u603_o;
  wire _al_u604_o;
  wire _al_u605_o;
  wire _al_u607_o;
  wire _al_u608_o;
  wire _al_u609_o;
  wire _al_u610_o;
  wire _al_u611_o;
  wire _al_u612_o;
  wire _al_u613_o;
  wire _al_u614_o;
  wire _al_u615_o;
  wire _al_u616_o;
  wire _al_u617_o;
  wire _al_u618_o;
  wire _al_u619_o;
  wire _al_u620_o;
  wire _al_u621_o;
  wire _al_u622_o;
  wire _al_u623_o;
  wire _al_u624_o;
  wire _al_u625_o;
  wire _al_u626_o;
  wire _al_u628_o;
  wire _al_u629_o;
  wire _al_u630_o;
  wire _al_u631_o;
  wire _al_u632_o;
  wire _al_u633_o;
  wire _al_u634_o;
  wire _al_u635_o;
  wire _al_u636_o;
  wire _al_u637_o;
  wire _al_u638_o;
  wire _al_u639_o;
  wire _al_u640_o;
  wire _al_u641_o;
  wire _al_u642_o;
  wire _al_u643_o;
  wire _al_u644_o;
  wire _al_u645_o;
  wire _al_u646_o;
  wire _al_u647_o;
  wire _al_u649_o;
  wire _al_u650_o;
  wire _al_u651_o;
  wire _al_u652_o;
  wire _al_u653_o;
  wire _al_u654_o;
  wire _al_u655_o;
  wire _al_u656_o;
  wire _al_u657_o;
  wire _al_u658_o;
  wire _al_u659_o;
  wire _al_u660_o;
  wire _al_u661_o;
  wire _al_u662_o;
  wire _al_u663_o;
  wire _al_u664_o;
  wire _al_u665_o;
  wire _al_u666_o;
  wire _al_u667_o;
  wire _al_u668_o;
  wire _al_u670_o;
  wire _al_u671_o;
  wire _al_u672_o;
  wire _al_u673_o;
  wire _al_u674_o;
  wire _al_u675_o;
  wire _al_u676_o;
  wire _al_u677_o;
  wire _al_u678_o;
  wire _al_u679_o;
  wire _al_u680_o;
  wire _al_u681_o;
  wire _al_u682_o;
  wire _al_u683_o;
  wire _al_u684_o;
  wire _al_u685_o;
  wire _al_u686_o;
  wire _al_u687_o;
  wire _al_u688_o;
  wire _al_u689_o;
  wire _al_u691_o;
  wire _al_u692_o;
  wire _al_u693_o;
  wire _al_u694_o;
  wire _al_u695_o;
  wire _al_u696_o;
  wire _al_u697_o;
  wire _al_u698_o;
  wire _al_u699_o;
  wire _al_u700_o;
  wire _al_u701_o;
  wire _al_u702_o;
  wire _al_u703_o;
  wire _al_u704_o;
  wire _al_u705_o;
  wire _al_u706_o;
  wire _al_u707_o;
  wire _al_u708_o;
  wire _al_u709_o;
  wire _al_u710_o;
  wire _al_u712_o;
  wire _al_u713_o;
  wire _al_u714_o;
  wire _al_u715_o;
  wire _al_u716_o;
  wire _al_u717_o;
  wire _al_u718_o;
  wire _al_u719_o;
  wire _al_u720_o;
  wire _al_u721_o;
  wire _al_u722_o;
  wire _al_u723_o;
  wire _al_u724_o;
  wire _al_u725_o;
  wire _al_u726_o;
  wire _al_u727_o;
  wire _al_u728_o;
  wire _al_u729_o;
  wire _al_u730_o;
  wire _al_u731_o;
  wire _al_u733_o;
  wire _al_u734_o;
  wire _al_u735_o;
  wire _al_u736_o;
  wire _al_u737_o;
  wire _al_u738_o;
  wire _al_u739_o;
  wire _al_u740_o;
  wire _al_u741_o;
  wire _al_u742_o;
  wire _al_u743_o;
  wire _al_u744_o;
  wire _al_u745_o;
  wire _al_u746_o;
  wire _al_u747_o;
  wire _al_u748_o;
  wire _al_u749_o;
  wire _al_u750_o;
  wire _al_u751_o;
  wire _al_u752_o;
  wire _al_u754_o;
  wire _al_u755_o;
  wire _al_u756_o;
  wire _al_u757_o;
  wire _al_u758_o;
  wire _al_u759_o;
  wire _al_u760_o;
  wire _al_u761_o;
  wire _al_u762_o;
  wire _al_u763_o;
  wire _al_u764_o;
  wire _al_u765_o;
  wire _al_u766_o;
  wire _al_u767_o;
  wire _al_u768_o;
  wire _al_u769_o;
  wire _al_u770_o;
  wire _al_u771_o;
  wire _al_u772_o;
  wire _al_u773_o;
  wire _al_u775_o;
  wire _al_u776_o;
  wire _al_u777_o;
  wire _al_u778_o;
  wire _al_u779_o;
  wire _al_u780_o;
  wire _al_u781_o;
  wire _al_u782_o;
  wire _al_u783_o;
  wire _al_u784_o;
  wire _al_u785_o;
  wire _al_u786_o;
  wire _al_u787_o;
  wire _al_u788_o;
  wire _al_u789_o;
  wire _al_u790_o;
  wire _al_u791_o;
  wire _al_u792_o;
  wire _al_u793_o;
  wire _al_u794_o;
  wire _al_u796_o;
  wire _al_u797_o;
  wire _al_u798_o;
  wire _al_u799_o;
  wire _al_u800_o;
  wire _al_u801_o;
  wire _al_u802_o;
  wire _al_u803_o;
  wire _al_u804_o;
  wire _al_u805_o;
  wire _al_u806_o;
  wire _al_u807_o;
  wire _al_u808_o;
  wire _al_u809_o;
  wire _al_u810_o;
  wire _al_u811_o;
  wire _al_u812_o;
  wire _al_u813_o;
  wire _al_u814_o;
  wire _al_u815_o;
  wire _al_u817_o;
  wire _al_u818_o;
  wire _al_u819_o;
  wire _al_u820_o;
  wire _al_u821_o;
  wire _al_u822_o;
  wire _al_u823_o;
  wire _al_u824_o;
  wire _al_u825_o;
  wire _al_u826_o;
  wire _al_u827_o;
  wire _al_u828_o;
  wire _al_u829_o;
  wire _al_u830_o;
  wire _al_u831_o;
  wire _al_u832_o;
  wire _al_u833_o;
  wire _al_u834_o;
  wire _al_u835_o;
  wire _al_u836_o;
  wire _al_u838_o;
  wire _al_u839_o;
  wire _al_u840_o;
  wire _al_u841_o;
  wire _al_u842_o;
  wire _al_u843_o;
  wire _al_u844_o;
  wire _al_u845_o;
  wire _al_u846_o;
  wire _al_u847_o;
  wire _al_u848_o;
  wire _al_u849_o;
  wire _al_u850_o;
  wire _al_u851_o;
  wire _al_u852_o;
  wire _al_u853_o;
  wire _al_u854_o;
  wire _al_u855_o;
  wire _al_u856_o;
  wire _al_u857_o;
  wire _al_u859_o;
  wire _al_u860_o;
  wire _al_u861_o;
  wire _al_u862_o;
  wire _al_u863_o;
  wire _al_u864_o;
  wire _al_u865_o;
  wire _al_u866_o;
  wire _al_u867_o;
  wire _al_u868_o;
  wire _al_u869_o;
  wire _al_u870_o;
  wire _al_u871_o;
  wire _al_u872_o;
  wire _al_u873_o;
  wire _al_u874_o;
  wire _al_u875_o;
  wire _al_u876_o;
  wire _al_u877_o;
  wire _al_u878_o;
  wire _al_u880_o;
  wire _al_u881_o;
  wire _al_u882_o;
  wire _al_u883_o;
  wire _al_u884_o;
  wire _al_u885_o;
  wire _al_u886_o;
  wire _al_u887_o;
  wire _al_u888_o;
  wire _al_u889_o;
  wire _al_u890_o;
  wire _al_u891_o;
  wire _al_u892_o;
  wire _al_u893_o;
  wire _al_u894_o;
  wire _al_u895_o;
  wire _al_u896_o;
  wire _al_u897_o;
  wire _al_u898_o;
  wire _al_u899_o;
  wire _al_u901_o;
  wire _al_u902_o;
  wire _al_u903_o;
  wire _al_u904_o;
  wire _al_u905_o;
  wire _al_u906_o;
  wire _al_u907_o;
  wire _al_u908_o;
  wire _al_u909_o;
  wire _al_u910_o;
  wire _al_u911_o;
  wire _al_u912_o;
  wire _al_u913_o;
  wire _al_u914_o;
  wire _al_u915_o;
  wire _al_u916_o;
  wire _al_u917_o;
  wire _al_u918_o;
  wire _al_u919_o;
  wire _al_u920_o;
  wire _al_u922_o;
  wire _al_u923_o;
  wire _al_u924_o;
  wire _al_u925_o;
  wire _al_u926_o;
  wire _al_u927_o;
  wire _al_u928_o;
  wire _al_u929_o;
  wire _al_u930_o;
  wire _al_u931_o;
  wire _al_u932_o;
  wire _al_u933_o;
  wire _al_u934_o;
  wire _al_u935_o;
  wire _al_u936_o;
  wire _al_u937_o;
  wire _al_u938_o;
  wire _al_u939_o;
  wire _al_u940_o;
  wire _al_u941_o;
  wire _al_u943_o;
  wire _al_u944_o;
  wire _al_u945_o;
  wire _al_u946_o;
  wire _al_u947_o;
  wire _al_u948_o;
  wire _al_u949_o;
  wire _al_u950_o;
  wire _al_u951_o;
  wire _al_u952_o;
  wire _al_u953_o;
  wire _al_u954_o;
  wire _al_u955_o;
  wire _al_u956_o;
  wire _al_u957_o;
  wire _al_u958_o;
  wire _al_u959_o;
  wire _al_u960_o;
  wire _al_u961_o;
  wire _al_u962_o;
  wire _al_u964_o;
  wire _al_u965_o;
  wire _al_u966_o;
  wire _al_u967_o;
  wire _al_u968_o;
  wire _al_u969_o;
  wire _al_u970_o;
  wire _al_u971_o;
  wire _al_u972_o;
  wire _al_u973_o;
  wire _al_u974_o;
  wire _al_u975_o;
  wire _al_u976_o;
  wire _al_u977_o;
  wire _al_u978_o;
  wire _al_u979_o;
  wire _al_u980_o;
  wire _al_u981_o;
  wire _al_u982_o;
  wire _al_u983_o;
  wire _al_u985_o;
  wire _al_u986_o;
  wire _al_u987_o;
  wire _al_u988_o;
  wire _al_u989_o;
  wire _al_u990_o;
  wire _al_u991_o;
  wire _al_u992_o;
  wire _al_u993_o;
  wire _al_u994_o;
  wire _al_u995_o;
  wire _al_u996_o;
  wire _al_u997_o;
  wire _al_u998_o;
  wire _al_u999_o;
  wire \cfg_int/wrapper_cfg_inst/rst ;  // D:/td/td/cw\cfg_int.v(23)
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_1 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_13 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_15 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ;
  wire \cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ;
  wire \cfg_int/wrapper_cfg_inst/shift_0 ;  // D:/td/td/cw\cfg_int.v(23)
  wire \cfg_int/wrapper_cfg_inst/tap_inst/jscan_1_r ;  // D:/td/td/cw\tap.v(16)
  wire \cfg_int/wrapper_cfg_inst/tap_inst/jscan_1_r2 ;  // D:/td/td/cw\tap.v(17)
  wire clock_pad;  // __top.v(4)
  wire control_0;
  wire control_1;
  wire control_10;
  wire control_100;
  wire control_101;
  wire control_102;
  wire control_103;
  wire control_104;
  wire control_105;
  wire control_106;
  wire control_107;
  wire control_108;
  wire control_109;
  wire control_11;
  wire control_110;
  wire control_111;
  wire control_112;
  wire control_113;
  wire control_114;
  wire control_115;
  wire control_116;
  wire control_117;
  wire control_118;
  wire control_119;
  wire control_12;
  wire control_120;
  wire control_121;
  wire control_122;
  wire control_123;
  wire control_124;
  wire control_125;
  wire control_126;
  wire control_127;
  wire control_128;
  wire control_129;
  wire control_13;
  wire control_130;
  wire control_131;
  wire control_132;
  wire control_133;
  wire control_134;
  wire control_135;
  wire control_136;
  wire control_137;
  wire control_138;
  wire control_139;
  wire control_14;
  wire control_140;
  wire control_141;
  wire control_142;
  wire control_143;
  wire control_144;
  wire control_145;
  wire control_146;
  wire control_147;
  wire control_148;
  wire control_149;
  wire control_15;
  wire control_150;
  wire control_151;
  wire control_152;
  wire control_153;
  wire control_154;
  wire control_155;
  wire control_156;
  wire control_157;
  wire control_158;
  wire control_159;
  wire control_16;
  wire control_160;
  wire control_161;
  wire control_162;
  wire control_163;
  wire control_164;
  wire control_165;
  wire control_166;
  wire control_167;
  wire control_168;
  wire control_169;
  wire control_17;
  wire control_170;
  wire control_171;
  wire control_172;
  wire control_173;
  wire control_174;
  wire control_175;
  wire control_176;
  wire control_177;
  wire control_178;
  wire control_179;
  wire control_18;
  wire control_180;
  wire control_181;
  wire control_182;
  wire control_183;
  wire control_184;
  wire control_185;
  wire control_186;
  wire control_187;
  wire control_188;
  wire control_189;
  wire control_19;
  wire control_190;
  wire control_191;
  wire control_192;
  wire control_193;
  wire control_194;
  wire control_195;
  wire control_196;
  wire control_197;
  wire control_198;
  wire control_199;
  wire control_2;
  wire control_20;
  wire control_200;
  wire control_201;
  wire control_202;
  wire control_203;
  wire control_204;
  wire control_205;
  wire control_206;
  wire control_207;
  wire control_208;
  wire control_209;
  wire control_21;
  wire control_210;
  wire control_211;
  wire control_212;
  wire control_213;
  wire control_214;
  wire control_215;
  wire control_216;
  wire control_217;
  wire control_218;
  wire control_219;
  wire control_22;
  wire control_220;
  wire control_221;
  wire control_222;
  wire control_223;
  wire control_224;
  wire control_225;
  wire control_226;
  wire control_227;
  wire control_228;
  wire control_229;
  wire control_23;
  wire control_230;
  wire control_231;
  wire control_232;
  wire control_233;
  wire control_234;
  wire control_235;
  wire control_236;
  wire control_237;
  wire control_238;
  wire control_239;
  wire control_24;
  wire control_240;
  wire control_241;
  wire control_242;
  wire control_243;
  wire control_244;
  wire control_245;
  wire control_246;
  wire control_247;
  wire control_248;
  wire control_249;
  wire control_25;
  wire control_250;
  wire control_251;
  wire control_252;
  wire control_253;
  wire control_254;
  wire control_255;
  wire control_256;
  wire control_257;
  wire control_258;
  wire control_259;
  wire control_26;
  wire control_260;
  wire control_261;
  wire control_262;
  wire control_263;
  wire control_264;
  wire control_265;
  wire control_266;
  wire control_267;
  wire control_268;
  wire control_269;
  wire control_27;
  wire control_270;
  wire control_271;
  wire control_272;
  wire control_273;
  wire control_274;
  wire control_275;
  wire control_276;
  wire control_277;
  wire control_278;
  wire control_279;
  wire control_28;
  wire control_280;
  wire control_281;
  wire control_282;
  wire control_283;
  wire control_284;
  wire control_285;
  wire control_286;
  wire control_287;
  wire control_288;
  wire control_289;
  wire control_29;
  wire control_290;
  wire control_291;
  wire control_292;
  wire control_293;
  wire control_294;
  wire control_295;
  wire control_296;
  wire control_297;
  wire control_298;
  wire control_299;
  wire control_3;
  wire control_30;
  wire control_300;
  wire control_301;
  wire control_302;
  wire control_303;
  wire control_304;
  wire control_305;
  wire control_306;
  wire control_307;
  wire control_308;
  wire control_309;
  wire control_31;
  wire control_310;
  wire control_311;
  wire control_312;
  wire control_32;
  wire control_33;
  wire control_34;
  wire control_35;
  wire control_36;
  wire control_37;
  wire control_38;
  wire control_39;
  wire control_40;
  wire control_41;
  wire control_42;
  wire control_43;
  wire control_44;
  wire control_45;
  wire control_46;
  wire control_47;
  wire control_48;
  wire control_49;
  wire control_50;
  wire control_51;
  wire control_52;
  wire control_53;
  wire control_54;
  wire control_55;
  wire control_56;
  wire control_57;
  wire control_58;
  wire control_59;
  wire control_6;
  wire control_60;
  wire control_61;
  wire control_62;
  wire control_63;
  wire control_64;
  wire control_65;
  wire control_66;
  wire control_67;
  wire control_68;
  wire control_69;
  wire control_7;
  wire control_70;
  wire control_71;
  wire control_72;
  wire control_73;
  wire control_74;
  wire control_75;
  wire control_76;
  wire control_77;
  wire control_78;
  wire control_79;
  wire control_8;
  wire control_80;
  wire control_81;
  wire control_82;
  wire control_83;
  wire control_84;
  wire control_85;
  wire control_86;
  wire control_87;
  wire control_88;
  wire control_89;
  wire control_9;
  wire control_90;
  wire control_91;
  wire control_92;
  wire control_93;
  wire control_94;
  wire control_95;
  wire control_96;
  wire control_97;
  wire control_98;
  wire control_99;
  wire jrstn;
  wire jscan_0;
  wire jscan_1;
  wire jshift;
  wire jtck;
  wire jtck_leading;
  wire jtdi;
  wire jtdo_0;
  wire jtdo_1;
  wire jupdate;
  wire lt0_c1;
  wire lt0_c11;
  wire lt0_c13;
  wire lt0_c15;
  wire lt0_c17;
  wire lt0_c19;
  wire lt0_c21;
  wire lt0_c23;
  wire lt0_c25;
  wire lt0_c27;
  wire lt0_c29;
  wire lt0_c3;
  wire lt0_c31;
  wire lt0_c5;
  wire lt0_c7;
  wire lt0_c9;
  wire \m/dram_c0_mode ;
  wire \m/dram_c0_wclk ;
  wire \m/dram_c0_we ;
  wire \m/dram_c1_mode ;
  wire \m/dram_c1_wclk ;
  wire \m/dram_c1_we ;
  wire \m/dram_c2_mode ;
  wire \m/dram_c2_wclk ;
  wire \m/dram_c2_we ;
  wire \m/dram_c3_mode ;
  wire \m/dram_c3_wclk ;
  wire \m/dram_c3_we ;
  wire \m/dram_c4_mode ;
  wire \m/dram_c4_wclk ;
  wire \m/dram_c4_we ;
  wire \m/dram_c5_mode ;
  wire \m/dram_c5_wclk ;
  wire \m/dram_c5_we ;
  wire \m/dram_c6_mode ;
  wire \m/dram_c6_wclk ;
  wire \m/dram_c6_we ;
  wire \m/dram_c7_mode ;
  wire \m/dram_c7_wclk ;
  wire \m/dram_c7_we ;
  wire memwrite_cs;  // __top.v(14)
  wire n0;
  wire n7;
  wire rst_pad;  // __top.v(3)
  wire status_0;
  wire status_1;
  wire status_10;
  wire status_11;
  wire status_12;
  wire status_13;
  wire status_14;
  wire status_15;
  wire status_16;
  wire status_17;
  wire status_2;
  wire status_3;
  wire status_4;
  wire status_5;
  wire status_6;
  wire status_7;
  wire status_8;
  wire status_9;
  wire \t/a/EX_operation$0$_lutinv_placeOpt_1 ;
  wire \t/a/EX_operation$0$_lutinv_placeOpt_2 ;
  wire \t/a/EX_operation$0$_lutinv_placeOpt_3 ;
  wire \t/a/EX_operation$0$_lutinv_placeOpt_4 ;
  wire \t/a/EX_operation$0$_lutinv_placeOpt_5 ;
  wire \t/a/ID_rs1$0$_placeOpt_1 ;
  wire \t/a/ID_rs1$0$_placeOpt_10 ;
  wire \t/a/ID_rs1$0$_placeOpt_11 ;
  wire \t/a/ID_rs1$0$_placeOpt_12 ;
  wire \t/a/ID_rs1$0$_placeOpt_13 ;
  wire \t/a/ID_rs1$0$_placeOpt_14 ;
  wire \t/a/ID_rs1$0$_placeOpt_15 ;
  wire \t/a/ID_rs1$0$_placeOpt_16 ;
  wire \t/a/ID_rs1$0$_placeOpt_17 ;
  wire \t/a/ID_rs1$0$_placeOpt_18 ;
  wire \t/a/ID_rs1$0$_placeOpt_19 ;
  wire \t/a/ID_rs1$0$_placeOpt_2 ;
  wire \t/a/ID_rs1$0$_placeOpt_20 ;
  wire \t/a/ID_rs1$0$_placeOpt_21 ;
  wire \t/a/ID_rs1$0$_placeOpt_3 ;
  wire \t/a/ID_rs1$0$_placeOpt_4 ;
  wire \t/a/ID_rs1$0$_placeOpt_5 ;
  wire \t/a/ID_rs1$0$_placeOpt_6 ;
  wire \t/a/ID_rs1$0$_placeOpt_7 ;
  wire \t/a/ID_rs1$0$_placeOpt_8 ;
  wire \t/a/ID_rs1$0$_placeOpt_9 ;
  wire \t/a/ID_rs1$1$_placeOpt_1 ;
  wire \t/a/ID_rs1$1$_placeOpt_10 ;
  wire \t/a/ID_rs1$1$_placeOpt_11 ;
  wire \t/a/ID_rs1$1$_placeOpt_12 ;
  wire \t/a/ID_rs1$1$_placeOpt_13 ;
  wire \t/a/ID_rs1$1$_placeOpt_14 ;
  wire \t/a/ID_rs1$1$_placeOpt_15 ;
  wire \t/a/ID_rs1$1$_placeOpt_16 ;
  wire \t/a/ID_rs1$1$_placeOpt_17 ;
  wire \t/a/ID_rs1$1$_placeOpt_18 ;
  wire \t/a/ID_rs1$1$_placeOpt_19 ;
  wire \t/a/ID_rs1$1$_placeOpt_2 ;
  wire \t/a/ID_rs1$1$_placeOpt_20 ;
  wire \t/a/ID_rs1$1$_placeOpt_21 ;
  wire \t/a/ID_rs1$1$_placeOpt_3 ;
  wire \t/a/ID_rs1$1$_placeOpt_4 ;
  wire \t/a/ID_rs1$1$_placeOpt_5 ;
  wire \t/a/ID_rs1$1$_placeOpt_6 ;
  wire \t/a/ID_rs1$1$_placeOpt_7 ;
  wire \t/a/ID_rs1$1$_placeOpt_8 ;
  wire \t/a/ID_rs1$1$_placeOpt_9 ;
  wire \t/a/ID_rs1$2$_placeOpt_1 ;
  wire \t/a/ID_rs1$2$_placeOpt_10 ;
  wire \t/a/ID_rs1$2$_placeOpt_2 ;
  wire \t/a/ID_rs1$2$_placeOpt_3 ;
  wire \t/a/ID_rs1$2$_placeOpt_4 ;
  wire \t/a/ID_rs1$2$_placeOpt_5 ;
  wire \t/a/ID_rs1$2$_placeOpt_6 ;
  wire \t/a/ID_rs1$2$_placeOpt_7 ;
  wire \t/a/ID_rs1$2$_placeOpt_8 ;
  wire \t/a/ID_rs1$2$_placeOpt_9 ;
  wire \t/a/ID_rs1$3$_placeOpt_1 ;
  wire \t/a/ID_rs1$3$_placeOpt_2 ;
  wire \t/a/ID_rs1$3$_placeOpt_3 ;
  wire \t/a/ID_rs2$0$_placeOpt_1 ;
  wire \t/a/ID_rs2$0$_placeOpt_10 ;
  wire \t/a/ID_rs2$0$_placeOpt_11 ;
  wire \t/a/ID_rs2$0$_placeOpt_12 ;
  wire \t/a/ID_rs2$0$_placeOpt_13 ;
  wire \t/a/ID_rs2$0$_placeOpt_14 ;
  wire \t/a/ID_rs2$0$_placeOpt_15 ;
  wire \t/a/ID_rs2$0$_placeOpt_16 ;
  wire \t/a/ID_rs2$0$_placeOpt_17 ;
  wire \t/a/ID_rs2$0$_placeOpt_18 ;
  wire \t/a/ID_rs2$0$_placeOpt_19 ;
  wire \t/a/ID_rs2$0$_placeOpt_2 ;
  wire \t/a/ID_rs2$0$_placeOpt_20 ;
  wire \t/a/ID_rs2$0$_placeOpt_21 ;
  wire \t/a/ID_rs2$0$_placeOpt_22 ;
  wire \t/a/ID_rs2$0$_placeOpt_3 ;
  wire \t/a/ID_rs2$0$_placeOpt_4 ;
  wire \t/a/ID_rs2$0$_placeOpt_5 ;
  wire \t/a/ID_rs2$0$_placeOpt_6 ;
  wire \t/a/ID_rs2$0$_placeOpt_7 ;
  wire \t/a/ID_rs2$0$_placeOpt_8 ;
  wire \t/a/ID_rs2$0$_placeOpt_9 ;
  wire \t/a/ID_rs2$1$_placeOpt_1 ;
  wire \t/a/ID_rs2$1$_placeOpt_10 ;
  wire \t/a/ID_rs2$1$_placeOpt_11 ;
  wire \t/a/ID_rs2$1$_placeOpt_12 ;
  wire \t/a/ID_rs2$1$_placeOpt_13 ;
  wire \t/a/ID_rs2$1$_placeOpt_14 ;
  wire \t/a/ID_rs2$1$_placeOpt_15 ;
  wire \t/a/ID_rs2$1$_placeOpt_16 ;
  wire \t/a/ID_rs2$1$_placeOpt_17 ;
  wire \t/a/ID_rs2$1$_placeOpt_18 ;
  wire \t/a/ID_rs2$1$_placeOpt_19 ;
  wire \t/a/ID_rs2$1$_placeOpt_2 ;
  wire \t/a/ID_rs2$1$_placeOpt_20 ;
  wire \t/a/ID_rs2$1$_placeOpt_21 ;
  wire \t/a/ID_rs2$1$_placeOpt_3 ;
  wire \t/a/ID_rs2$1$_placeOpt_4 ;
  wire \t/a/ID_rs2$1$_placeOpt_5 ;
  wire \t/a/ID_rs2$1$_placeOpt_6 ;
  wire \t/a/ID_rs2$1$_placeOpt_7 ;
  wire \t/a/ID_rs2$1$_placeOpt_8 ;
  wire \t/a/ID_rs2$1$_placeOpt_9 ;
  wire \t/a/ID_rs2$2$_placeOpt_1 ;
  wire \t/a/ID_rs2$2$_placeOpt_10 ;
  wire \t/a/ID_rs2$2$_placeOpt_2 ;
  wire \t/a/ID_rs2$2$_placeOpt_3 ;
  wire \t/a/ID_rs2$2$_placeOpt_4 ;
  wire \t/a/ID_rs2$2$_placeOpt_5 ;
  wire \t/a/ID_rs2$2$_placeOpt_6 ;
  wire \t/a/ID_rs2$2$_placeOpt_7 ;
  wire \t/a/ID_rs2$2$_placeOpt_8 ;
  wire \t/a/ID_rs2$2$_placeOpt_9 ;
  wire \t/a/ID_rs2$3$_placeOpt_1 ;
  wire \t/a/ID_rs2$3$_placeOpt_2 ;
  wire \t/a/ID_rs2$3$_placeOpt_3 ;
  wire \t/a/WB_regwritecs ;  // cpu.v(69)
  wire \t/a/alu/add0/c11 ;
  wire \t/a/alu/add0/c15 ;
  wire \t/a/alu/add0/c19 ;
  wire \t/a/alu/add0/c23 ;
  wire \t/a/alu/add0/c27 ;
  wire \t/a/alu/add0/c3 ;
  wire \t/a/alu/add0/c31 ;
  wire \t/a/alu/add0/c7 ;
  wire \t/a/alu/lt0_c1 ;
  wire \t/a/alu/lt0_c11 ;
  wire \t/a/alu/lt0_c13 ;
  wire \t/a/alu/lt0_c15 ;
  wire \t/a/alu/lt0_c17 ;
  wire \t/a/alu/lt0_c19 ;
  wire \t/a/alu/lt0_c21 ;
  wire \t/a/alu/lt0_c23 ;
  wire \t/a/alu/lt0_c25 ;
  wire \t/a/alu/lt0_c27 ;
  wire \t/a/alu/lt0_c29 ;
  wire \t/a/alu/lt0_c3 ;
  wire \t/a/alu/lt0_c31 ;
  wire \t/a/alu/lt0_c5 ;
  wire \t/a/alu/lt0_c7 ;
  wire \t/a/alu/lt0_c9 ;
  wire \t/a/alu/n104_lutinv ;
  wire \t/a/alu/n105_lutinv ;
  wire \t/a/alu/n106_lutinv ;
  wire \t/a/alu/n132_lutinv ;
  wire \t/a/alu/n133_lutinv ;
  wire \t/a/alu/n134_lutinv ;
  wire \t/a/alu/n135_lutinv ;
  wire \t/a/alu/n136_lutinv ;
  wire \t/a/alu/n137_lutinv ;
  wire \t/a/alu/n138_lutinv ;
  wire \t/a/alu/n142_lutinv ;
  wire \t/a/alu/n143_lutinv ;
  wire \t/a/alu/n144_lutinv ;
  wire \t/a/alu/n145_lutinv ;
  wire \t/a/alu/n146_lutinv ;
  wire \t/a/alu/n147_lutinv ;
  wire \t/a/alu/n148_lutinv ;
  wire \t/a/alu/n149_lutinv ;
  wire \t/a/alu/n150_lutinv ;
  wire \t/a/alu/n151_lutinv ;
  wire \t/a/alu/n152_lutinv ;
  wire \t/a/alu/n153_lutinv ;
  wire \t/a/alu/n154_lutinv ;
  wire \t/a/alu/n155_lutinv ;
  wire \t/a/alu/n156_lutinv ;
  wire \t/a/alu/n157_lutinv ;
  wire \t/a/alu/n158_lutinv ;
  wire \t/a/alu/n159_lutinv ;
  wire \t/a/alu/n160_lutinv ;
  wire \t/a/alu/n161_lutinv ;
  wire \t/a/alu/n162_lutinv ;
  wire \t/a/alu/n163_lutinv ;
  wire \t/a/alu/n164_lutinv ;
  wire \t/a/alu/n165_lutinv ;
  wire \t/a/alu/n166_lutinv ;
  wire \t/a/alu/n167_lutinv ;
  wire \t/a/alu/n168_lutinv ;
  wire \t/a/alu/n169_lutinv ;
  wire \t/a/alu/n170_lutinv ;
  wire \t/a/alu/n173_lutinv ;
  wire \t/a/alu/n17_lutinv ;
  wire \t/a/alu/n18_lutinv ;
  wire \t/a/alu/n19_lutinv ;
  wire \t/a/alu/n202_lutinv ;
  wire \t/a/alu/n204_lutinv ;
  wire \t/a/alu/n20_lutinv ;
  wire \t/a/alu/n21_lutinv ;
  wire \t/a/alu/n22_lutinv ;
  wire \t/a/alu/n232_lutinv ;
  wire \t/a/alu/n233_lutinv ;
  wire \t/a/alu/n234_lutinv ;
  wire \t/a/alu/n23_lutinv ;
  wire \t/a/alu/n24_lutinv ;
  wire \t/a/alu/n25_lutinv ;
  wire \t/a/alu/n260_lutinv ;
  wire \t/a/alu/n261_lutinv ;
  wire \t/a/alu/n262_lutinv ;
  wire \t/a/alu/n263_lutinv ;
  wire \t/a/alu/n264_lutinv ;
  wire \t/a/alu/n265_lutinv ;
  wire \t/a/alu/n266_lutinv ;
  wire \t/a/alu/n26_lutinv ;
  wire \t/a/alu/n27_lutinv ;
  wire \t/a/alu/n28_lutinv ;
  wire \t/a/alu/n29_lutinv ;
  wire \t/a/alu/n30_lutinv ;
  wire \t/a/alu/n31_lutinv ;
  wire \t/a/alu/n32_lutinv ;
  wire \t/a/alu/n33_lutinv ;
  wire \t/a/alu/n34_lutinv ;
  wire \t/a/alu/n35_lutinv ;
  wire \t/a/alu/n36_lutinv ;
  wire \t/a/alu/n37_lutinv ;
  wire \t/a/alu/n38_lutinv ;
  wire \t/a/alu/n39_lutinv ;
  wire \t/a/alu/n40_lutinv ;
  wire \t/a/alu/n41_lutinv ;
  wire \t/a/alu/n42_lutinv ;
  wire \t/a/alu/n43_lutinv ;
  wire \t/a/alu/n44_lutinv ;
  wire \t/a/alu/n45_lutinv ;
  wire \t/a/alu/n56_lutinv ;
  wire \t/a/alu/n57_lutinv ;
  wire \t/a/alu/n8 ;
  wire \t/a/alu/sub0/c11 ;
  wire \t/a/alu/sub0/c15 ;
  wire \t/a/alu/sub0/c19 ;
  wire \t/a/alu/sub0/c23 ;
  wire \t/a/alu/sub0/c27 ;
  wire \t/a/alu/sub0/c3 ;
  wire \t/a/alu/sub0/c31 ;
  wire \t/a/alu/sub0/c7 ;
  wire \t/a/aluin/n10_lutinv ;
  wire \t/a/aluin/n11_lutinv ;
  wire \t/a/aluin/n12_lutinv ;
  wire \t/a/aluin/n35_lutinv ;
  wire \t/a/aluin/n5_lutinv ;
  wire \t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_1 ;
  wire \t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 ;
  wire \t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_3 ;
  wire \t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 ;
  wire \t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/condition/add0/c11 ;
  wire \t/a/condition/add0/c15 ;
  wire \t/a/condition/add0/c19 ;
  wire \t/a/condition/add0/c23 ;
  wire \t/a/condition/add0/c27 ;
  wire \t/a/condition/add0/c3 ;
  wire \t/a/condition/add0/c31 ;
  wire \t/a/condition/add0/c7 ;
  wire \t/a/condition/lt0_c1 ;
  wire \t/a/condition/lt0_c11 ;
  wire \t/a/condition/lt0_c13 ;
  wire \t/a/condition/lt0_c15 ;
  wire \t/a/condition/lt0_c17 ;
  wire \t/a/condition/lt0_c19 ;
  wire \t/a/condition/lt0_c21 ;
  wire \t/a/condition/lt0_c23 ;
  wire \t/a/condition/lt0_c25 ;
  wire \t/a/condition/lt0_c27 ;
  wire \t/a/condition/lt0_c29 ;
  wire \t/a/condition/lt0_c3 ;
  wire \t/a/condition/lt0_c31 ;
  wire \t/a/condition/lt0_c5 ;
  wire \t/a/condition/lt0_c7 ;
  wire \t/a/condition/lt0_c9 ;
  wire \t/a/condition/lt1_c1 ;
  wire \t/a/condition/lt1_c11 ;
  wire \t/a/condition/lt1_c13 ;
  wire \t/a/condition/lt1_c15 ;
  wire \t/a/condition/lt1_c17 ;
  wire \t/a/condition/lt1_c19 ;
  wire \t/a/condition/lt1_c21 ;
  wire \t/a/condition/lt1_c23 ;
  wire \t/a/condition/lt1_c25 ;
  wire \t/a/condition/lt1_c27 ;
  wire \t/a/condition/lt1_c29 ;
  wire \t/a/condition/lt1_c3 ;
  wire \t/a/condition/lt1_c31 ;
  wire \t/a/condition/lt1_c5 ;
  wire \t/a/condition/lt1_c7 ;
  wire \t/a/condition/lt1_c9 ;
  wire \t/a/condition/n0_lutinv ;
  wire \t/a/condition/n10 ;
  wire \t/a/condition/n1_lutinv ;
  wire \t/a/condition/n9 ;
  wire \t/a/ex_mem/n0 ;
  wire \t/a/if_id/n9 ;
  wire \t/a/instr/add0/c11 ;
  wire \t/a/instr/add0/c15 ;
  wire \t/a/instr/add0/c19 ;
  wire \t/a/instr/add0/c23 ;
  wire \t/a/instr/add0/c27 ;
  wire \t/a/instr/add0/c3 ;
  wire \t/a/instr/add0/c31 ;
  wire \t/a/instr/add0/c7 ;
  wire \t/a/instr/add2/c11 ;
  wire \t/a/instr/add2/c15 ;
  wire \t/a/instr/add2/c19 ;
  wire \t/a/instr/add2/c23 ;
  wire \t/a/instr/add2/c27 ;
  wire \t/a/instr/add2/c3 ;
  wire \t/a/instr/add2/c7 ;
  wire \t/a/n0_lutinv ;
  wire \t/a/n19 ;
  wire \t/a/n2 ;
  wire \t/a/n24_lutinv ;
  wire \t/a/n29 ;
  wire \t/a/n4_lutinv ;
  wire \t/a/n9_lutinv ;
  wire \t/a/regfile/mux39_b0_sel_is_3_o ;
  wire \t/a/regfile/mux39_b1000_sel_is_3_o ;
  wire \t/a/regfile/mux39_b100_sel_is_3_o ;
  wire \t/a/regfile/mux39_b128_sel_is_3_o ;
  wire \t/a/regfile/mux39_b160_sel_is_3_o ;
  wire \t/a/regfile/mux39_b192_sel_is_3_o ;
  wire \t/a/regfile/mux39_b224_sel_is_3_o ;
  wire \t/a/regfile/mux39_b256_sel_is_3_o ;
  wire \t/a/regfile/mux39_b288_sel_is_3_o ;
  wire \t/a/regfile/mux39_b320_sel_is_3_o ;
  wire \t/a/regfile/mux39_b32_sel_is_3_o ;
  wire \t/a/regfile/mux39_b352_sel_is_3_o ;
  wire \t/a/regfile/mux39_b384_sel_is_3_o ;
  wire \t/a/regfile/mux39_b416_sel_is_3_o ;
  wire \t/a/regfile/mux39_b448_sel_is_3_o ;
  wire \t/a/regfile/mux39_b480_sel_is_3_o ;
  wire \t/a/regfile/mux39_b512_sel_is_3_o ;
  wire \t/a/regfile/mux39_b544_sel_is_3_o ;
  wire \t/a/regfile/mux39_b576_sel_is_3_o ;
  wire \t/a/regfile/mux39_b608_sel_is_3_o ;
  wire \t/a/regfile/mux39_b640_sel_is_3_o ;
  wire \t/a/regfile/mux39_b64_sel_is_3_o ;
  wire \t/a/regfile/mux39_b672_sel_is_3_o ;
  wire \t/a/regfile/mux39_b704_sel_is_3_o ;
  wire \t/a/regfile/mux39_b736_sel_is_3_o ;
  wire \t/a/regfile/mux39_b768_sel_is_3_o ;
  wire \t/a/regfile/mux39_b800_sel_is_3_o ;
  wire \t/a/regfile/mux39_b832_sel_is_3_o ;
  wire \t/a/regfile/mux39_b864_sel_is_3_o ;
  wire \t/a/regfile/mux39_b896_sel_is_3_o ;
  wire \t/a/regfile/mux39_b928_sel_is_3_o ;
  wire \t/a/regfile/mux39_b960_sel_is_3_o ;
  wire \t/a/regfile/n1_lutinv ;
  wire \t/a/regfile/n3_lutinv ;
  wire \t/a/risk_jump/n11_lutinv ;
  wire \t/a/risk_jump/n19 ;
  wire \t/a/risk_jump/n24_lutinv ;
  wire \t/a/risk_jump/n35_lutinv ;
  wire \t/a/risk_jump/n42_lutinv ;
  wire \t/a/unconditional/eq1/or_xor_i0$5$_i1$5$_o_o_lutinv ;
  wire \t/busarbitration/mux5_b0_sel_is_3_o ;
  wire \t/busarbitration/mux6_b16_sel_is_3_o ;
  wire \t/busarbitration/n3 ;
  wire \t/busarbitration/n3_placeOpt_1 ;
  wire \t/busarbitration/n3_placeOpt_2 ;
  wire \t/busarbitration/n3_placeOpt_3 ;
  wire \t/busarbitration/n3_placeOpt_4 ;
  wire \t/busarbitration/n3_placeOpt_5 ;
  wire \t/instrnop ;  // top2.v(12)
  wire \t/instruction$2$_neg_lutinv ;
  wire \t/instruction$3$_neg_lutinv ;
  wire \t/instruction$4$_neg_lutinv ;
  wire \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r ;  // D:/td/td/cw\detecEdge.v(19)
  wire \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 ;
  wire \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 ;
  wire \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 ;
  wire \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 ;
  wire \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this ;  // D:/td/td/cw\detecEdge.v(17)
  wire \trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r ;  // D:/td/td/cw\detecEdge.v(18)
  wire \trig_node/trigger_node_int_0/add0/c1 ;
  wire \trig_node/trigger_node_int_0/add0/c11 ;
  wire \trig_node/trigger_node_int_0/add0/c13 ;
  wire \trig_node/trigger_node_int_0/add0/c3 ;
  wire \trig_node/trigger_node_int_0/add0/c5 ;
  wire \trig_node/trigger_node_int_0/add0/c7 ;
  wire \trig_node/trigger_node_int_0/add0/c9 ;
  wire \trig_node/trigger_node_int_0/add1/c11 ;
  wire \trig_node/trigger_node_int_0/add1/c15 ;
  wire \trig_node/trigger_node_int_0/add1/c3 ;
  wire \trig_node/trigger_node_int_0/add1/c7 ;
  wire \trig_node/trigger_node_int_0/emb_store_en ;  // D:/td/td/cw\trigger_node.v(75)
  wire \trig_node/trigger_node_int_0/force_acq_fin ;  // D:/td/td/cw\trigger_node.v(40)
  wire \trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ;
  wire \trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 ;
  wire \trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 ;
  wire \trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 ;
  wire \trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 ;
  wire \trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 ;
  wire \trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 ;
  wire \trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 ;
  wire \trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c11 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c15 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c3 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c7 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c11 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c15 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c3 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c7 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c1 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c11 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c13 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c15 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c3 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c5 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c7 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c9 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13$0$_en ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n19 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n2 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c11 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c15 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c3 ;
  wire \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c7 ;
  wire \trig_node/trigger_node_int_0/lt0_c1 ;
  wire \trig_node/trigger_node_int_0/lt0_c11 ;
  wire \trig_node/trigger_node_int_0/lt0_c13 ;
  wire \trig_node/trigger_node_int_0/lt0_c15 ;
  wire \trig_node/trigger_node_int_0/lt0_c3 ;
  wire \trig_node/trigger_node_int_0/lt0_c5 ;
  wire \trig_node/trigger_node_int_0/lt0_c7 ;
  wire \trig_node/trigger_node_int_0/lt0_c9 ;
  wire \trig_node/trigger_node_int_0/n177 ;
  wire \trig_node/trigger_node_int_0/pause_sync ;  // D:/td/td/cw\trigger_node.v(85)
  wire \trig_node/trigger_node_int_0/pause_sync0 ;  // D:/td/td/cw\trigger_node.v(85)
  wire \trig_node/trigger_node_int_0/sub0/c1 ;
  wire \trig_node/trigger_node_int_0/sub0/c11 ;
  wire \trig_node/trigger_node_int_0/sub0/c13 ;
  wire \trig_node/trigger_node_int_0/sub0/c15 ;
  wire \trig_node/trigger_node_int_0/sub0/c3 ;
  wire \trig_node/trigger_node_int_0/sub0/c5 ;
  wire \trig_node/trigger_node_int_0/sub0/c7 ;
  wire \trig_node/trigger_node_int_0/sub0/c9 ;
  wire \trig_node/trigger_node_int_0/trig_rstn_sync ;  // D:/td/td/cw\trigger_node.v(35)
  wire \trig_node/trigger_node_int_0/trig_rstn_sync0 ;  // D:/td/td/cw\trigger_node.v(35)
  wire \trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ;
  wire \trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ;
  wire \trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ;
  wire \trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ;
  wire \trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ;
  wire \trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ;
  wire \trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ;
  wire \trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ;
  wire \trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ;
  wire \trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ;
  wire \u1/c1 ;
  wire \u1/c11 ;
  wire \u1/c13 ;
  wire \u1/c15 ;
  wire \u1/c17 ;
  wire \u1/c19 ;
  wire \u1/c21 ;
  wire \u1/c23 ;
  wire \u1/c25 ;
  wire \u1/c27 ;
  wire \u1/c29 ;
  wire \u1/c3 ;
  wire \u1/c5 ;
  wire \u1/c7 ;
  wire \u1/c9 ;
  wire \u3/c11 ;
  wire \u3/c15 ;
  wire \u3/c19 ;
  wire \u3/c23 ;
  wire \u3/c27 ;
  wire \u3/c3 ;
  wire \u3/c7 ;
  wire wt_ce;

  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUT1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUT0(16'b0111000000110000),
    .INIT_LUT1(16'b1111000010110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1000 (
    .a({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/ID_rs1$0$_placeOpt_16 }),
    .b({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/ID_rs1$1$_placeOpt_16 }),
    .c({\t/a/ID_rs1$2$_placeOpt_6 ,\t/a/ID_rs1$2$_placeOpt_6 }),
    .d({\t/a/regfile/regfile$30$ [0],\t/a/regfile/regfile$30$ [0]}),
    .mi({open_n12,\t/a/regfile/regfile$31$ [0]}),
    .fx({open_n17,_al_u1000_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*B*A)"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(1*D*~C*B*A)"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1001|t/a/regfile/reg0_b928  (
    .a({_al_u1000_o,_al_u256_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_10 ,\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs1$1$_placeOpt_10 ,\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$28$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$29$ [0],\t/a/WB_rd [3]}),
    .mi({open_n21,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1001_o,\t/a/regfile/mux39_b928_sel_is_3_o }),
    .q({open_n36,\t/a/regfile/regfile$29$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1002|_al_u1718  (
    .a({\t/a/ID_rs1$0$_placeOpt_10 ,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/ID_rs1$1$_placeOpt_10 ,\t/a/ID_rs2$1$_placeOpt_12 }),
    .c({\t/a/ID_rs1$2$_placeOpt_4 ,\t/a/ID_rs2$2$_placeOpt_5 }),
    .d({\t/a/regfile/regfile$26$ [0],\t/a/regfile/regfile$26$ [0]}),
    .e({\t/a/regfile/regfile$27$ [0],\t/a/regfile/regfile$27$ [0]}),
    .f({_al_u1002_o,_al_u1718_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(C*~((~A*~B))*~(D)+C*(~A*~B)*~(D)+~(C)*(~A*~B)*D+C*(~A*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(C*~((~A*~B))*~(D)+C*(~A*~B)*~(D)+~(C)*(~A*~B)*D+C*(~A*~B)*D))"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0001000111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1004|_al_u1003  (
    .a({_al_u1003_o,_al_u1002_o}),
    .b({_al_u1001_o,\t/a/ID_rs1$0$_placeOpt_10 }),
    .c({_al_u999_o,\t/a/ID_rs1$1$_placeOpt_10 }),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$24$ [0]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$25$ [0]}),
    .f({_al_u1004_o,_al_u1003_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*~(D*C))"),
    //.LUTF1("A*D*~B*~C+A*D*~B*C"),
    //.LUTG0("(~1*B*A*~(D*C))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0010001000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1006|_al_u1038  (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_fun3 [0],\t/a/MEM_regdat2 [0]}),
    .c({open_n81,\t/a/MEM_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .e({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [2]}),
    .mi({o_data[0],o_data[0]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({\t/busarbitration/mux6_b16_sel_is_3_o ,o_data[0]}),
    .q({\trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*A)"),
    //.LUT1("(B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010000010100000),
    .INIT_LUT1(16'b1100000011000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1007|_al_u1022  (
    .a({open_n98,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .b({\t/a/MEM_regdat2 [31],open_n99}),
    .c({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/a/MEM_regdat2 [16]}),
    .clk(clock_pad),
    .mi({o_data[16],o_data[16]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({o_data[31],o_data[16]}),
    .q({\trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*A)"),
    //.LUTF1("(C*A)"),
    //.LUTG0("(B*A)"),
    //.LUTG1("(C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b1010000010100000),
    .INIT_LUTG0(16'b1000100010001000),
    .INIT_LUTG1(16'b1010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1008|_al_u1021  (
    .a({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .b({open_n116,\t/a/MEM_regdat2 [17]}),
    .c({\t/a/MEM_regdat2 [30],open_n117}),
    .clk(clock_pad),
    .mi({o_data[17],o_data[17]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({o_data[30],o_data[17]}),
    .q({\trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1111000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1009|_al_u1020  (
    .c({\t/a/MEM_regdat2 [29],open_n142}),
    .clk(clock_pad),
    .d({open_n144,\t/a/MEM_regdat2 [18]}),
    .e({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .mi({o_data[29],o_data[29]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({o_data[29],o_data[18]}),
    .q({\trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*A)"),
    //.LUT1("(D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1010101000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1010|_al_u1019  (
    .a({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .b({open_n160,\t/a/MEM_regdat2 [19]}),
    .clk(clock_pad),
    .d({\t/a/MEM_regdat2 [28],open_n164}),
    .mi({o_data[28],o_data[28]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({o_data[28],o_data[19]}),
    .q({\trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*A)"),
    //.LUT1("(C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101000000000),
    .INIT_LUT1(16'b1010000010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1011|_al_u1018  (
    .a({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .c({\t/a/MEM_regdat2 [27],open_n180}),
    .clk(clock_pad),
    .d({open_n182,\t/a/MEM_regdat2 [20]}),
    .mi({o_data[27],o_data[27]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({o_data[27],o_data[20]}),
    .q({\trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*B)"),
    //.LUTF1("(C*B)"),
    //.LUTG0("(D*B)"),
    //.LUTG1("(C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110000000000),
    .INIT_LUTF1(16'b1100000011000000),
    .INIT_LUTG0(16'b1100110000000000),
    .INIT_LUTG1(16'b1100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1012|_al_u1017  (
    .b({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .c({\t/a/MEM_regdat2 [26],open_n198}),
    .clk(clock_pad),
    .d({open_n200,\t/a/MEM_regdat2 [21]}),
    .mi({o_data[26],o_data[26]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({o_data[26],o_data[21]}),
    .q({\trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("0"),
    //.LUTG0("(C*D)"),
    //.LUTG1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1013|_al_u1016  (
    .c({open_n222,\t/a/MEM_regdat2 [22]}),
    .clk(clock_pad),
    .d({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .e({\t/a/MEM_regdat2 [25],open_n224}),
    .mi({o_data[25],o_data[25]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({o_data[25],o_data[22]}),
    .q({\trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*A)"),
    //.LUT1("(B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010000010100000),
    .INIT_LUT1(16'b1000100010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1014|_al_u1015  (
    .a({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .b({\t/a/MEM_regdat2 [24],open_n240}),
    .c({open_n241,\t/a/MEM_regdat2 [23]}),
    .clk(clock_pad),
    .mi({o_data[24],o_data[24]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f(o_data[24:23]),
    .q({\trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*~(D*C))"),
    //.LUTF1("(~0*B*C*(A@D))"),
    //.LUTG0("(~1*B*A*~(D*C))"),
    //.LUTG1("(~1*B*C*(A@D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0100000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1023|_al_u1035  (
    .a({\t/a/MEM_fun3 [1],memwrite_cs}),
    .b({\t/a/MEM_regdat2 [9],\t/a/MEM_regdat2 [3]}),
    .c({memwrite_cs,\t/a/MEM_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [1]}),
    .e({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [2]}),
    .mi({o_data[9],o_data[9]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({o_data[9],o_data[3]}),
    .q({\trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*~(D*C))"),
    //.LUTF1("(~0*C*A*(B@D))"),
    //.LUTG0("(~1*B*A*~(D*C))"),
    //.LUTG1("(~1*C*A*(B@D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0010000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1024|_al_u1034  (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_fun3 [1],\t/a/MEM_regdat2 [4]}),
    .c({\t/a/MEM_regdat2 [8],\t/a/MEM_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [1]}),
    .e({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [2]}),
    .mi({o_data[8],o_data[8]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({o_data[8],o_data[4]}),
    .q({\trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*~(D*C))"),
    //.LUTF1("(~0*B*C*(A@D))"),
    //.LUTG0("(~1*B*A*~(D*C))"),
    //.LUTG1("(~1*B*C*(A@D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0100000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1025|_al_u1031  (
    .a({\t/a/MEM_fun3 [1],memwrite_cs}),
    .b({\t/a/MEM_regdat2 [15],\t/a/MEM_regdat2 [7]}),
    .c({memwrite_cs,\t/a/MEM_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [1]}),
    .e({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [2]}),
    .mi({o_data[15],o_data[15]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({o_data[15],o_data[7]}),
    .q({\trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*(D@C))"),
    //.LUTF1("(~0*C*A*(B@D))"),
    //.LUTG0("(~1*B*A*(D@C))"),
    //.LUTG1("(~1*C*A*(B@D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100010000000),
    .INIT_LUTF1(16'b0010000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1026|_al_u1030  (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_fun3 [1],\t/a/MEM_regdat2 [10]}),
    .c({\t/a/MEM_regdat2 [14],\t/a/MEM_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [1]}),
    .e({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [2]}),
    .mi({o_data[14],o_data[14]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .f({o_data[14],o_data[10]}),
    .q({\trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*(D@C))"),
    //.LUT1("(~1*B*A*(C@D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100010000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    _al_u1028 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [12],\t/a/MEM_regdat2 [12]}),
    .c(\t/a/MEM_fun3 [1:0]),
    .clk(clock_pad),
    .d({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [1]}),
    .mi({o_data[12],\t/a/MEM_fun3 [2]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .fx({open_n336,o_data[12]}),
    .q({\trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/level_0_r ,open_n337}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*(D@C))"),
    //.LUT1("(~1*B*A*(D@C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100010000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    _al_u1029 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [11],\t/a/MEM_regdat2 [11]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .mi({o_data[11],\t/a/MEM_fun3 [2]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .fx({open_n352,o_data[11]}),
    .q({\trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/level_0_r ,open_n353}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*~(D*C))"),
    //.LUT1("(~1*B*A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    _al_u1032 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [6],\t/a/MEM_regdat2 [6]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .mi({o_data[6],\t/a/MEM_fun3 [2]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .fx({open_n368,o_data[6]}),
    .q({\trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/level_0_r ,open_n369}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*~(D*C))"),
    //.LUT1("(~1*B*A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    _al_u1033 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [5],\t/a/MEM_regdat2 [5]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .mi({o_data[5],\t/a/MEM_fun3 [2]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .fx({open_n384,o_data[5]}),
    .q({\trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/level_0_r ,open_n385}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*~(D*C))"),
    //.LUT1("(~1*B*A*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    _al_u1036 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [2],\t/a/MEM_regdat2 [2]}),
    .c(\t/a/MEM_fun3 [1:0]),
    .clk(clock_pad),
    .d({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [1]}),
    .mi({o_data[2],\t/a/MEM_fun3 [2]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .fx({open_n400,o_data[2]}),
    .q({\trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/level_0_r ,open_n401}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*~(D*C))"),
    //.LUT1("(~1*B*A*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    _al_u1037 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [1],\t/a/MEM_regdat2 [1]}),
    .c(\t/a/MEM_fun3 [1:0]),
    .clk(clock_pad),
    .d({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [1]}),
    .mi({o_data[1],\t/a/MEM_fun3 [2]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .fx({open_n416,o_data[1]}),
    .q({\trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/level_0_r ,open_n417}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000010101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1039|t/a/if_id/reg5_b5  (
    .a({addr[5],open_n418}),
    .b({open_n419,\t/a/MEM_aludat [5]}),
    .c({open_n420,\t/memstraddress [5]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({memwrite_cs,\t/busarbitration/n3_placeOpt_5 }),
    .mi({open_n431,\t/memstraddress [5]}),
    .sr(rst_pad),
    .f({n3[3],addr[5]}),
    .q({open_n435,\t/a/ID_memstraddr [5]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    //.LUT1("(~D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101011001100),
    .INIT_LUT1(16'b0000000010101010),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1040|_al_u297  (
    .a({addr[4],\t/memstraddress [4]}),
    .b({open_n436,\t/a/MEM_aludat [4]}),
    .clk(clock_pad),
    .d({memwrite_cs,\t/busarbitration/n3_placeOpt_5 }),
    .mi({addr[4],addr[4]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({n3[2],addr[4]}),
    .q({\trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000010101010),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1041|_al_u300  (
    .a({addr[3],open_n453}),
    .b({open_n454,\t/a/MEM_aludat [3]}),
    .c({open_n455,\t/memstraddress [3]}),
    .clk(clock_pad),
    .d({memwrite_cs,\t/busarbitration/n3_placeOpt_3 }),
    .mi({addr[3],addr[3]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .f({n3[1],addr[3]}),
    .q({\trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*D*~C*~A+B*D*~C*~A+~B*D*C*~A+B*D*C*~A"),
    //.LUTF1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~B*D*~C*~A+B*D*~C*~A+~B*D*C*~A+B*D*C*~A+~B*~D*~C*A+B*~D*~C*A+~B*D*~C*A+B*D*~C*A+~B*~D*C*A+B*~D*C*A+~B*D*C*A+B*D*C*A"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010100000000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b1111111110101010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1042|_al_u311  (
    .a({open_n470,\t/busarbitration/n3_placeOpt_4 }),
    .clk(clock_pad),
    .d({addr[2],\t/a/MEM_aludat [2]}),
    .e({memwrite_cs,\t/memstraddress [2]}),
    .mi({addr[2],addr[2]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .f({n3[0],addr[2]}),
    .q({\trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0@C)*~(D*~B))"),
    //.LUT1("(~A*~(1@C)*~(D*~B))"),
    .INIT_LUT0(16'b0000010000000101),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1044 (
    .a({_al_u1043_o,_al_u1043_o}),
    .b({\t/a/ID_rs2$2$_placeOpt_7 ,\t/a/ID_rs2$2$_placeOpt_7 }),
    .c({\t/a/ID_rs2 [4],\t/a/ID_rs2 [4]}),
    .d({\t/a/WB_rd [2],\t/a/WB_rd [2]}),
    .mi({open_n503,\t/a/WB_rd [4]}),
    .fx({open_n508,_al_u1044_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~0*C)*~(D*~B))"),
    //.LUT1("(A*~(~1*D)*~(C*~B))"),
    .INIT_LUT0(16'b0000100000001010),
    .INIT_LUT1(16'b1000101010001010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1045 (
    .a({_al_u1044_o,_al_u1044_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/ID_rs2$0$_placeOpt_21 }),
    .c({\t/a/WB_rd [0],\t/a/ID_rs2$2$_placeOpt_7 }),
    .d({\t/a/ID_rs2$2$_placeOpt_7 ,\t/a/WB_rd [0]}),
    .mi({open_n523,\t/a/WB_rd [2]}),
    .fx({open_n528,_al_u1045_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(A*B)"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(A*B)"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1048|_al_u1047  (
    .a({_al_u1047_o,_al_u1046_o}),
    .b({_al_u1045_o,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({open_n531,\t/a/ID_rs2$3$_placeOpt_3 }),
    .d({open_n534,\t/a/WB_rd [1]}),
    .e({open_n535,\t/a/WB_rd [3]}),
    .f({\t/a/regfile/n3_lutinv ,_al_u1047_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*~B*A)"),
    //.LUTF1("(B*D)"),
    //.LUTG0("(1*D*~C*~B*A)"),
    //.LUTG1("(B*D)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1100110000000000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b1100110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1049|_al_u2604  (
    .a({open_n556,\t/a/regfile/n3_lutinv }),
    .b({\t/a/WB_regwritecs ,\t/a/risk_jump/n42_lutinv }),
    .c({open_n557,\t/a/risk_jump/n35_lutinv }),
    .d({\t/a/regfile/n3_lutinv ,\t/a/n19 }),
    .e({open_n560,\t/a/condition/n1_lutinv }),
    .f({_al_u1049_o,_al_u2604_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("A*~B*~C*~D+A*~B*C*~D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0001000100110011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1050|_al_u1505  (
    .a({\t/a/ID_rs2$0$_placeOpt_8 ,_al_u1501_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_16 ,_al_u1502_o}),
    .c({open_n581,_al_u1503_o}),
    .d({\t/a/regfile/regfile$5$ [9],_al_u1504_o}),
    .e({\t/a/regfile/regfile$4$ [9],\t/a/ID_rs2$2$_placeOpt_8 }),
    .f({_al_u1050_o,_al_u1505_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1053|t/a/regfile/reg0_b73  (
    .a({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/regfile/regfile$2$ [9]}),
    .b({\t/a/ID_rs2$1$_placeOpt_11 ,\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/regfile/regfile$3$ [9],\t/a/regfile/regfile$3$ [9]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [9],\t/a/ID_rs1$0$_placeOpt_10 }),
    .mi({open_n614,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u1053_o,_al_u347_o}),
    .q({open_n618,\t/a/regfile/regfile$2$ [9]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1054 (
    .a({_al_u1050_o,_al_u1050_o}),
    .b({_al_u1051_o,_al_u1051_o}),
    .c({_al_u1052_o,_al_u1052_o}),
    .d({_al_u1053_o,_al_u1053_o}),
    .mi({open_n631,\t/a/ID_rs2$2$_placeOpt_10 }),
    .fx({open_n636,_al_u1054_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1059|t/a/regfile/reg0_b425  (
    .a({_al_u1056_o,_al_u1055_o}),
    .b({_al_u1054_o,\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1058_o,\t/a/regfile/regfile$12$ [9]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [9]}),
    .mi({open_n640,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u1059_o,_al_u1056_o}),
    .q({open_n655,\t/a/regfile/regfile$13$ [9]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1064 (
    .a({_al_u1060_o,_al_u1060_o}),
    .b({_al_u1061_o,_al_u1061_o}),
    .c({_al_u1062_o,_al_u1062_o}),
    .d({_al_u1063_o,_al_u1063_o}),
    .mi({open_n668,\t/a/ID_rs2$2$_placeOpt_1 }),
    .fx({open_n673,_al_u1064_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1069|t/a/regfile/reg0_b937  (
    .a({_al_u1064_o,_al_u1065_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_16 }),
    .c({_al_u1068_o,\t/a/ID_rs2$1$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1066_o,\t/a/regfile/regfile$28$ [9]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [9]}),
    .mi({open_n677,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u1069_o,_al_u1066_o}),
    .q({open_n692,\t/a/regfile/regfile$29$ [9]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~A*B*~D*~C+A*B*~D*~C+A*B*D*~C+~A*B*~D*C"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*B*~D*~C+A*B*~D*~C+A*B*D*~C+~A*B*~D*C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1072|t/a/regfile/reg0_b968  (
    .a({\t/a/ID_rs2$0$_placeOpt_16 ,\t/a/regfile/regfile$30$ [8]}),
    .b({\t/a/ID_rs2$1$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$31$ [8],\t/a/ID_rs1$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [8],\t/a/regfile/regfile$31$ [8]}),
    .e({open_n693,\t/a/ID_rs1$0$_placeOpt_2 }),
    .mi({open_n695,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u1072_o,_al_u370_o}),
    .q({open_n710,\t/a/regfile/regfile$30$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1075|_al_u1285  (
    .a({_al_u1071_o,_al_u1281_o}),
    .b({_al_u1072_o,_al_u1282_o}),
    .c({_al_u1073_o,_al_u1283_o}),
    .d({_al_u1074_o,_al_u1284_o}),
    .e({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/ID_rs2$2$_placeOpt_1 }),
    .f({_al_u1075_o,_al_u1285_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100000011000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1080|t/a/regfile/reg0_b680  (
    .a({_al_u1077_o,_al_u1076_o}),
    .b({_al_u1075_o,\t/a/ID_rs2$0$_placeOpt_6 }),
    .c({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1079_o,\t/a/regfile/regfile$20$ [8]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [8]}),
    .mi({open_n734,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u1080_o,_al_u1077_o}),
    .q({open_n749,\t/a/regfile/regfile$21$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+D*~B*C*A"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~D*~B*~C*~A+~D*~B*~C*A"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1081|_al_u1327  (
    .a({open_n750,_al_u1323_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_19 ,_al_u1324_o}),
    .c({\t/a/regfile/regfile$4$ [8],_al_u1325_o}),
    .d({\t/a/ID_rs2$0$_placeOpt_14 ,_al_u1326_o}),
    .e({\t/a/regfile/regfile$5$ [8],\t/a/ID_rs2$2$_placeOpt_6 }),
    .f({_al_u1081_o,_al_u1327_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1082|_al_u1369  (
    .a({\t/a/ID_rs2$0$_placeOpt_3 ,_al_u1365_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_13 ,_al_u1366_o}),
    .c({\t/a/regfile/regfile$6$ [8],_al_u1367_o}),
    .d({\t/a/regfile/regfile$7$ [8],_al_u1368_o}),
    .e({open_n775,\t/a/ID_rs2$2$_placeOpt_6 }),
    .f({_al_u1082_o,_al_u1369_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1084|t/a/regfile/reg0_b72  (
    .a({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/regfile/regfile$2$ [8]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1$1$_placeOpt_13 }),
    .c({\t/a/regfile/regfile$3$ [8],\t/a/regfile/regfile$3$ [8]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [8],\t/a/ID_rs1$0$_placeOpt_10 }),
    .mi({open_n806,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u1084_o,_al_u358_o}),
    .q({open_n810,\t/a/regfile/regfile$2$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011011100000100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1090|t/a/regfile/reg0_b424  (
    .a({_al_u1087_o,_al_u1086_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_20 }),
    .c({_al_u1089_o,\t/a/ID_rs2$1$_placeOpt_18 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1085_o,\t/a/regfile/regfile$12$ [8]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [8]}),
    .mi({open_n812,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u1090_o,_al_u1087_o}),
    .q({open_n827,\t/a/regfile/regfile$13$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~A*~C)*~((~B*~D))*~(0)+(~A*~C)*(~B*~D)*~(0)+~((~A*~C))*(~B*~D)*0+(~A*~C)*(~B*~D)*0)"),
    //.LUTF1("~D*~B*~A*~C+D*~B*~A*~C+D*~B*A*~C+~D*~B*~A*C+D*~B*~A*C+D*~B*A*C"),
    //.LUTG0("~((~A*~C)*~((~B*~D))*~(1)+(~A*~C)*(~B*~D)*~(1)+~((~A*~C))*(~B*~D)*1+(~A*~C)*(~B*~D)*1)"),
    //.LUTG1("~D*~B*~A*~C+~D*~B*~A*C"),
    .INIT_LUTF0(16'b1111101011111010),
    .INIT_LUTF1(16'b0011001100010001),
    .INIT_LUTG0(16'b1111111111001100),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1092|_al_u1096  (
    .a({\t/a/regfile/regfile$4$ [7],_al_u1095_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_13 ,_al_u1093_o}),
    .c({open_n828,_al_u1094_o}),
    .d({\t/a/ID_rs2$0$_placeOpt_3 ,_al_u1092_o}),
    .e({\t/a/regfile/regfile$5$ [7],\t/a/ID_rs2$2$_placeOpt_6 }),
    .f({_al_u1092_o,_al_u1096_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1095|t/a/regfile/reg0_b71  (
    .a({\t/a/ID_rs2 [0],\t/a/regfile/regfile$2$ [7]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1$1$_placeOpt_13 }),
    .c({\t/a/regfile/regfile$3$ [7],\t/a/regfile/regfile$3$ [7]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [7],\t/a/ID_rs1$0$_placeOpt_13 }),
    .mi({open_n861,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({_al_u1095_o,_al_u389_o}),
    .q({open_n865,\t/a/regfile/regfile$2$ [7]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1101|t/a/regfile/reg0_b423  (
    .a({_al_u1096_o,_al_u1097_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_10 }),
    .c({_al_u1100_o,\t/a/ID_rs2$1$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1098_o,\t/a/regfile/regfile$12$ [7]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [7]}),
    .mi({open_n867,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({_al_u1101_o,_al_u1098_o}),
    .q({open_n882,\t/a/regfile/regfile$13$ [7]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1106|_al_u1421  (
    .a({_al_u1102_o,_al_u1417_o}),
    .b({_al_u1103_o,_al_u1418_o}),
    .c({_al_u1104_o,_al_u1419_o}),
    .d({_al_u1105_o,_al_u1420_o}),
    .e({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/ID_rs2$2$_placeOpt_1 }),
    .f({_al_u1106_o,_al_u1421_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1111|t/a/regfile/reg0_b935  (
    .a({_al_u1108_o,_al_u1107_o}),
    .b({_al_u1106_o,\t/a/ID_rs2$0$_placeOpt_16 }),
    .c({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1110_o,\t/a/regfile/regfile$28$ [7]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [7]}),
    .mi({open_n906,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({_al_u1111_o,_al_u1108_o}),
    .q({open_n921,\t/a/regfile/regfile$29$ [7]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1113|t/a/regfile/reg0_b134  (
    .a({\t/a/regfile/regfile$4$ [6],_al_u2606_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_21 ,_al_u2610_o}),
    .c({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/MEM_aludat [6]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [6],\t/a/reg_writedat [6]}),
    .mi({open_n932,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u1113_o,_al_u2730_o}),
    .q({open_n936,\t/a/regfile/regfile$4$ [6]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100000101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1116|t/a/regfile/reg0_b70  (
    .a({\t/a/ID_rs2$1$_placeOpt_18 ,\t/a/regfile/regfile$2$ [6]}),
    .b({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs1$1$_placeOpt_18 }),
    .c({\t/a/regfile/regfile$3$ [6],\t/a/regfile/regfile$3$ [6]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [6],\t/a/ID_rs1$0$_placeOpt_18 }),
    .mi({open_n947,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u1116_o,_al_u400_o}),
    .q({open_n951,\t/a/regfile/regfile$2$ [6]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1117 (
    .a({_al_u1113_o,_al_u1113_o}),
    .b({_al_u1114_o,_al_u1114_o}),
    .c({_al_u1115_o,_al_u1115_o}),
    .d({_al_u1116_o,_al_u1116_o}),
    .mi({open_n964,\t/a/ID_rs2$2$_placeOpt_4 }),
    .fx({open_n969,_al_u1117_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1122|t/a/regfile/reg0_b422  (
    .a({_al_u1117_o,_al_u1118_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_9 }),
    .c({_al_u1121_o,\t/a/ID_rs2$1$_placeOpt_17 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1119_o,\t/a/regfile/regfile$12$ [6]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [6]}),
    .mi({open_n973,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u1122_o,_al_u1119_o}),
    .q({open_n988,\t/a/regfile/regfile$13$ [6]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1127 (
    .a({_al_u1123_o,_al_u1123_o}),
    .b({_al_u1124_o,_al_u1124_o}),
    .c({_al_u1125_o,_al_u1125_o}),
    .d({_al_u1126_o,_al_u1126_o}),
    .mi({open_n1001,\t/a/ID_rs2$2$_placeOpt_2 }),
    .fx({open_n1006,_al_u1127_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1132|t/a/regfile/reg0_b934  (
    .a({_al_u1129_o,_al_u1128_o}),
    .b({_al_u1127_o,\t/a/ID_rs2$0$_placeOpt_19 }),
    .c({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_19 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1131_o,\t/a/regfile/regfile$28$ [6]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [6]}),
    .mi({open_n1010,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u1132_o,_al_u1129_o}),
    .q({open_n1025,\t/a/regfile/regfile$29$ [6]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1134|t/a/regfile/reg0_b133  (
    .a({\t/a/ID_rs2$0$_placeOpt_22 ,_al_u2606_o_placeOpt_2}),
    .b({\t/a/ID_rs2$1$_placeOpt_11 ,_al_u2610_o_placeOpt_2}),
    .c({\t/a/regfile/regfile$4$ [5],\t/a/MEM_aludat [5]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [5],\t/a/reg_writedat [5]}),
    .mi({open_n1036,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u1134_o,_al_u2737_o}),
    .q({open_n1040,\t/a/regfile/regfile$4$ [5]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~B*~C)*~((~D*~A))*~(0)+(~B*~C)*(~D*~A)*~(0)+~((~B*~C))*(~D*~A)*0+(~B*~C)*(~D*~A)*0)"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+~A*B*C*D"),
    //.LUTG0("~((~B*~C)*~((~D*~A))*~(1)+(~B*~C)*(~D*~A)*~(1)+~((~B*~C))*(~D*~A)*1+(~B*~C)*(~D*~A)*1)"),
    //.LUTG1("A*B*~C*~D+A*B*C*~D"),
    .INIT_LUTF0(16'b1111110011111100),
    .INIT_LUTF1(16'b0100010011001100),
    .INIT_LUTG0(16'b1111111110101010),
    .INIT_LUTG1(16'b0000000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1135|_al_u1138  (
    .a({\t/a/ID_rs2$0$_placeOpt_10 ,_al_u1134_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_11 ,_al_u1137_o}),
    .c({open_n1041,_al_u1136_o}),
    .d({\t/a/regfile/regfile$7$ [5],_al_u1135_o}),
    .e({\t/a/regfile/regfile$6$ [5],\t/a/ID_rs2$2$_placeOpt_10 }),
    .f({_al_u1135_o,_al_u1138_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1137|t/a/regfile/reg0_b69  (
    .a({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/regfile/regfile$2$ [5]}),
    .b({\t/a/ID_rs2$1$_placeOpt_12 ,\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/regfile/regfile$3$ [5],\t/a/regfile/regfile$3$ [5]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [5],\t/a/ID_rs1$0$_placeOpt_10 }),
    .mi({open_n1074,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u1137_o,_al_u421_o}),
    .q({open_n1078,\t/a/regfile/regfile$2$ [5]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1143|t/a/regfile/reg0_b421  (
    .a({_al_u1138_o,_al_u1139_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_9 }),
    .c({_al_u1142_o,\t/a/ID_rs2$1$_placeOpt_18 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1140_o,\t/a/regfile/regfile$12$ [5]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [5]}),
    .mi({open_n1080,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u1143_o,_al_u1140_o}),
    .q({open_n1095,\t/a/regfile/regfile$13$ [5]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1148|_al_u1358  (
    .a({_al_u1144_o,_al_u1354_o}),
    .b({_al_u1145_o,_al_u1355_o}),
    .c({_al_u1146_o,_al_u1356_o}),
    .d({_al_u1147_o,_al_u1357_o}),
    .e({\t/a/ID_rs2$2$_placeOpt_2 ,\t/a/ID_rs2$2$_placeOpt_2 }),
    .f({_al_u1148_o,_al_u1358_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1153|t/a/regfile/reg0_b933  (
    .a({_al_u1148_o,_al_u1149_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_18 }),
    .c({_al_u1152_o,\t/a/ID_rs2$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1150_o,\t/a/regfile/regfile$28$ [5]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [5]}),
    .mi({open_n1119,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u1153_o,_al_u1150_o}),
    .q({open_n1134,\t/a/regfile/regfile$29$ [5]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1155|t/a/regfile/reg0_b164  (
    .a({\t/a/regfile/regfile$5$ [4],_al_u2606_o_placeOpt_2}),
    .b({\t/a/regfile/regfile$4$ [4],_al_u2610_o_placeOpt_2}),
    .c({\t/a/ID_rs2$1$_placeOpt_11 ,\t/a/MEM_aludat [4]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/reg_writedat [4]}),
    .mi({open_n1145,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u1155_o,_al_u2742_o}),
    .q({open_n1149,\t/a/regfile/regfile$5$ [4]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~A*~(~0*B)))"),
    //.LUTF1("0"),
    //.LUTG0("~(C*~(D*~A*~(~1*B)))"),
    //.LUTG1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+B*~A*C*~D+B*A*C*~D+~B*~A*~C*D+~B*A*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0101111100001111),
    .INIT_LUTG1(16'b0000001111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1156|t/a/regfile/reg0_b196  (
    .a({open_n1150,_al_u1999_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$6$ [4],_al_u2000_o}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [4],\t/a/aluin/n10_lutinv }),
    .e({\t/a/ID_rs2$1$_placeOpt_11 ,\t/a/reg_writedat [4]}),
    .mi({open_n1152,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u1156_o,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .q({open_n1167,\t/a/regfile/regfile$6$ [4]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*C*B*A)"),
    //.LUTF1("~A*C*~D*~B+A*C*~D*~B+~A*C*D*~B+~A*C*~D*B+A*C*~D*B+~A*C*D*B"),
    //.LUTG0("(~1*~D*C*B*A)"),
    //.LUTG1("A*C*~D*~B+A*C*~D*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0101000011110000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1158|t/a/regfile/reg0_b100  (
    .a({\t/a/ID_rs2$0$_placeOpt_22 ,_al_u254_o}),
    .b({open_n1168,\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs2$1$_placeOpt_11 ,\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$3$ [4],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$2$ [4],\t/a/WB_rd [3]}),
    .mi({open_n1170,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u1158_o,\t/a/regfile/mux39_b100_sel_is_3_o }),
    .q({open_n1185,\t/a/regfile/regfile$3$ [4]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1164|t/a/regfile/reg0_b420  (
    .a({_al_u1161_o,_al_u1160_o}),
    .b({_al_u1159_o,\t/a/ID_rs2$0$_placeOpt_22 }),
    .c({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_12 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1163_o,\t/a/regfile/regfile$12$ [4]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [4]}),
    .mi({open_n1187,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u1164_o,_al_u1161_o}),
    .q({open_n1202,\t/a/regfile/regfile$13$ [4]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1169|_al_u1316  (
    .a({_al_u1165_o,_al_u1312_o}),
    .b({_al_u1166_o,_al_u1313_o}),
    .c({_al_u1167_o,_al_u1314_o}),
    .d({_al_u1168_o,_al_u1315_o}),
    .e({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/ID_rs2$2$_placeOpt_1 }),
    .f({_al_u1169_o,_al_u1316_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1174|t/a/regfile/reg0_b932  (
    .a({_al_u1169_o,_al_u1170_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_10 }),
    .c({_al_u1173_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1171_o,\t/a/regfile/regfile$28$ [4]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [4]}),
    .mi({open_n1226,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u1174_o,_al_u1171_o}),
    .q({open_n1241,\t/a/regfile/regfile$29$ [4]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1180|_al_u1222  (
    .a({_al_u1176_o,_al_u1218_o}),
    .b({_al_u1177_o,_al_u1219_o}),
    .c({_al_u1178_o,_al_u1220_o}),
    .d({_al_u1179_o,_al_u1221_o}),
    .e({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/ID_rs2$2$_placeOpt_1 }),
    .f({_al_u1180_o,_al_u1222_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1000100010001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1185|t/a/regfile/reg0_b675  (
    .a({_al_u1180_o,_al_u1181_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_16 }),
    .c({_al_u1184_o,\t/a/ID_rs2$1$_placeOpt_16 }),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1182_o,\t/a/regfile/regfile$20$ [3]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [3]}),
    .mi({open_n1265,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u1185_o,_al_u1182_o}),
    .q({open_n1280,\t/a/regfile/regfile$21$ [3]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000001100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1186|t/a/regfile/reg0_b131  (
    .a({\t/a/regfile/regfile$4$ [3],_al_u2614_o}),
    .b({\t/a/regfile/regfile$5$ [3],_al_u2616_o_placeOpt_3}),
    .c({\t/a/ID_rs2 [1],\t/a/MEM_aludat [3]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_10 ,\t/a/reg_writedat [3]}),
    .mi({open_n1291,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u1186_o,_al_u2752_o}),
    .q({open_n1295,\t/a/regfile/regfile$4$ [3]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~A*~(~0*B)))"),
    //.LUTF1("B*~A*~C*~D+B*A*~C*~D+B*~A*~C*D+B*A*~C*D"),
    //.LUTG0("~(C*~(D*~A*~(~1*B)))"),
    //.LUTG1("B*~A*~C*~D+B*A*~C*~D+B*~A*C*~D+B*A*C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0000110000001100),
    .INIT_LUTG0(16'b0101111100001111),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1187|t/a/regfile/reg0_b195  (
    .a({open_n1296,_al_u2009_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$6$ [3],_al_u2010_o}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [3],\t/a/aluin/n10_lutinv }),
    .e({\t/a/ID_rs2$0$_placeOpt_10 ,\t/a/reg_writedat [3]}),
    .mi({open_n1298,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u1187_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .q({open_n1313,\t/a/regfile/regfile$6$ [3]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~A*~(~0*B)))"),
    //.LUTF1("~D*B*~C*~A+D*B*~C*~A+~D*B*C*~A+~D*B*~C*A+D*B*~C*A+~D*B*C*A"),
    //.LUTG0("~(C*~(D*~A*~(~1*B)))"),
    //.LUTG1("D*B*~C*~A+D*B*~C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0101111100001111),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1187|t/a/regfile/reg0_b195_placeOpt_1  (
    .a({open_n1314,_al_u2009_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$7$ [3],_al_u2010_o}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_10 ,\t/a/aluin/n10_lutinv }),
    .e({\t/a/regfile/regfile$6$ [3],\t/a/reg_writedat [3]}),
    .mi({open_n1316,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({open_n1328,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_1 }));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~A*~(~0*B)))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*~C*D+A*B*~C*D"),
    //.LUTG0("~(C*~(D*~A*~(~1*B)))"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b0101111100001111),
    .INIT_LUTG1(16'b0000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1187|t/a/regfile/reg0_b195_placeOpt_2  (
    .a({\t/a/ID_rs2 [1],_al_u2009_o}),
    .b({open_n1334,\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$6$ [3],_al_u2010_o}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [3],\t/a/aluin/n10_lutinv }),
    .e({\t/a/ID_rs2$0$_placeOpt_10 ,\t/a/reg_writedat [3]}),
    .mi({open_n1336,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({open_n1348,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 }));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~A*~(~0*B)))"),
    //.LUTF1("D*~B*~A*~C+D*B*~A*~C+D*~B*A*~C+D*B*A*~C+D*~B*~A*C+D*~B*A*C"),
    //.LUTG0("~(C*~(D*~A*~(~1*B)))"),
    //.LUTG1("D*B*~A*~C+D*B*A*~C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0011111100000000),
    .INIT_LUTG0(16'b0101111100001111),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1187|t/a/regfile/reg0_b195_placeOpt_3  (
    .a({open_n1354,_al_u2009_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_10 ,\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$7$ [3],_al_u2010_o}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [1],\t/a/aluin/n10_lutinv }),
    .e({\t/a/regfile/regfile$6$ [3],\t/a/reg_writedat [3]}),
    .mi({open_n1356,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({open_n1368,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_3 }));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~A*~(~0*B)))"),
    //.LUTF1("0"),
    //.LUTG0("~(C*~(D*~A*~(~1*B)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*~B*~C*D+A*B*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0101111100001111),
    .INIT_LUTG1(16'b0000101001011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1187|t/a/regfile/reg0_b195_placeOpt_4  (
    .a({\t/a/ID_rs2$0$_placeOpt_10 ,_al_u2009_o}),
    .b({open_n1374,\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$7$ [3],_al_u2010_o}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$6$ [3],\t/a/aluin/n10_lutinv }),
    .e({\t/a/ID_rs2 [1],\t/a/reg_writedat [3]}),
    .mi({open_n1376,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({open_n1388,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1190 (
    .a({_al_u1186_o,_al_u1186_o}),
    .b({_al_u1187_o,_al_u1187_o}),
    .c({_al_u1188_o,_al_u1188_o}),
    .d({_al_u1189_o,_al_u1189_o}),
    .mi({open_n1406,\t/a/ID_rs2$2$_placeOpt_10 }),
    .fx({open_n1411,_al_u1190_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1195|t/a/regfile/reg0_b419  (
    .a({_al_u1192_o,_al_u1191_o}),
    .b({_al_u1190_o,\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1194_o,\t/a/regfile/regfile$12$ [3]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [3]}),
    .mi({open_n1415,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u1195_o,_al_u1192_o}),
    .q({open_n1430,\t/a/regfile/regfile$13$ [3]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*A*~C+~B*D*A*~C+~B*~D*A*C+~B*D*A*C"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D"),
    //.LUTG0("~B*~D*A*C+~B*D*A*C"),
    //.LUTG1("A*~B*~C*~D+A*~B*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000100010),
    .INIT_LUTF1(16'b0001001100010011),
    .INIT_LUTG0(16'b0010000000100000),
    .INIT_LUTG1(16'b0000001000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1197|t/a/regfile/reg0_b191  (
    .a({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/aluin/n5_lutinv }),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,_al_u1823_o}),
    .c({\t/a/regfile/regfile$5$ [31],\t/a/reg_writedat [31]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .e({\t/a/regfile/regfile$4$ [31],\t/a/alu_A_select [1]}),
    .mi({open_n1434,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1197_o,\t/a/aluin/sel0_b31/B0 }),
    .q({open_n1449,\t/a/regfile/regfile$5$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1200|t/a/regfile/reg0_b95  (
    .a({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/regfile/regfile$2$ [31]}),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/ID_rs1$1$_placeOpt_20 }),
    .c({\t/a/regfile/regfile$3$ [31],\t/a/regfile/regfile$3$ [31]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [31],\t/a/ID_rs1$0$_placeOpt_16 }),
    .mi({open_n1460,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1200_o,_al_u494_o}),
    .q({open_n1464,\t/a/regfile/regfile$2$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1201 (
    .a({_al_u1197_o,_al_u1197_o}),
    .b({_al_u1198_o,_al_u1198_o}),
    .c({_al_u1199_o,_al_u1199_o}),
    .d({_al_u1200_o,_al_u1200_o}),
    .mi({open_n1477,\t/a/ID_rs2$2$_placeOpt_7 }),
    .fx({open_n1482,_al_u1201_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000101000111010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1206|t/a/regfile/reg0_b447  (
    .a({_al_u1201_o,_al_u1202_o}),
    .b({_al_u1205_o,\t/a/ID_rs2$0$_placeOpt_21 }),
    .c({\t/a/ID_rs2$3$_placeOpt_3 ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1203_o,\t/a/regfile/regfile$12$ [31]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [31]}),
    .mi({open_n1486,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1206_o,_al_u1203_o}),
    .q({open_n1501,\t/a/regfile/regfile$13$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1211|_al_u1212  (
    .a({_al_u1207_o,\t/a/ID_rs2 [0]}),
    .b({_al_u1208_o,\t/a/ID_rs2 [1]}),
    .c({_al_u1209_o,\t/a/ID_rs2$2$_placeOpt_10 }),
    .d({_al_u1210_o,\t/a/regfile/regfile$31$ [31]}),
    .e({\t/a/ID_rs2$2$_placeOpt_10 ,\t/a/regfile/regfile$30$ [31]}),
    .f({_al_u1211_o,_al_u1212_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1216|t/a/regfile/reg0_b959  (
    .a({_al_u1211_o,_al_u1212_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_10 }),
    .c({_al_u1215_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1213_o,\t/a/regfile/regfile$28$ [31]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [31]}),
    .mi({open_n1525,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1216_o,_al_u1213_o}),
    .q({open_n1540,\t/a/regfile/regfile$29$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*~B*~C*D+A*B*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000101001011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1219|t/a/regfile/reg0_b990  (
    .a({\t/a/ID_rs2$0$_placeOpt_3 ,\t/a/regfile/regfile$30$ [30]}),
    .b({open_n1541,\t/a/ID_rs1$1$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$31$ [30],\t/a/ID_rs1$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [30],\t/a/regfile/regfile$31$ [30]}),
    .e({\t/a/ID_rs2$1$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_1 }),
    .mi({open_n1543,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1219_o,_al_u517_o}),
    .q({open_n1558,\t/a/regfile/regfile$30$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1000100010001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1227|t/a/regfile/reg0_b702  (
    .a({_al_u1222_o,_al_u1223_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_10 }),
    .c({_al_u1226_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1224_o,\t/a/regfile/regfile$20$ [30]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [30]}),
    .mi({open_n1560,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1227_o,_al_u1224_o}),
    .q({open_n1575,\t/a/regfile/regfile$21$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000010110101111),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1228|_al_u1232  (
    .a({\t/a/ID_rs2$0$_placeOpt_21 ,_al_u1228_o}),
    .b({open_n1576,_al_u1229_o}),
    .c({\t/a/regfile/regfile$4$ [30],_al_u1230_o}),
    .d({\t/a/regfile/regfile$5$ [30],_al_u1231_o}),
    .e({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/ID_rs2$2$_placeOpt_7 }),
    .f({_al_u1228_o,_al_u1232_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1231|t/a/regfile/reg0_b94  (
    .a({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/regfile/regfile$2$ [30]}),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/ID_rs1$1$_placeOpt_16 }),
    .c({\t/a/regfile/regfile$3$ [30],\t/a/regfile/regfile$3$ [30]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [30],\t/a/ID_rs1$0$_placeOpt_16 }),
    .mi({open_n1609,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1231_o,_al_u505_o}),
    .q({open_n1613,\t/a/regfile/regfile$2$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000010111001100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1237|t/a/regfile/reg0_b446  (
    .a({_al_u1234_o,_al_u1233_o}),
    .b({_al_u1232_o,\t/a/ID_rs2$0$_placeOpt_21 }),
    .c({_al_u1236_o,\t/a/ID_rs2$1$_placeOpt_15 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$3$_placeOpt_3 ,\t/a/regfile/regfile$12$ [30]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [30]}),
    .mi({open_n1615,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1237_o,_al_u1234_o}),
    .q({open_n1630,\t/a/regfile/regfile$13$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000000110101),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1239|t/a/regfile/reg0_b130  (
    .a({\t/a/regfile/regfile$4$ [2],_al_u2614_o}),
    .b({\t/a/regfile/regfile$5$ [2],_al_u2616_o}),
    .c({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/MEM_aludat [2]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_11 ,\t/a/reg_writedat [2]}),
    .mi({open_n1641,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u1239_o,_al_u2756_o}),
    .q({open_n1645,\t/a/regfile/regfile$4$ [2]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*(~A*~(0)*~(B)+~A*0*~(B)+~(~A)*0*B+~A*0*B)))"),
    //.LUTF1("~A*D*~B*~C+A*D*~B*~C+~A*D*B*~C+A*D*B*~C+~A*D*~B*C+~A*D*B*C"),
    //.LUTG0("~(C*~(D*(~A*~(1)*~(B)+~A*1*~(B)+~(~A)*1*B+~A*1*B)))"),
    //.LUTG1("A*D*~B*~C+A*D*B*~C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0101111100000000),
    .INIT_LUTG0(16'b1101111100001111),
    .INIT_LUTG1(16'b0000101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1240|t/a/regfile/reg0_b194  (
    .a({\t/a/ID_rs2$0$_placeOpt_21 ,_al_u2092_o}),
    .b({open_n1646,\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$7$ [2],_al_u2093_o}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/aluin/n10_lutinv }),
    .e({\t/a/regfile/regfile$6$ [2],\t/a/reg_writedat [2]}),
    .mi({open_n1648,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u1240_o,\t/a/EX_B [2]}),
    .q({open_n1663,\t/a/regfile/regfile$6$ [2]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1243 (
    .a({_al_u1239_o,_al_u1239_o}),
    .b({_al_u1240_o,_al_u1240_o}),
    .c({_al_u1241_o,_al_u1241_o}),
    .d({_al_u1242_o,_al_u1242_o}),
    .mi({open_n1676,\t/a/ID_rs2$2$_placeOpt_7 }),
    .fx({open_n1681,_al_u1243_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1248|t/a/regfile/reg0_b418  (
    .a({_al_u1243_o,_al_u1244_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_15 }),
    .c({_al_u1247_o,\t/a/ID_rs2$1$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1245_o,\t/a/regfile/regfile$12$ [2]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [2]}),
    .mi({open_n1685,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u1248_o,_al_u1245_o}),
    .q({open_n1700,\t/a/regfile/regfile$13$ [2]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111110110101000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1111110111111101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1253|_al_u1274  (
    .a({\t/a/ID_rs2 [2],_al_u1270_o}),
    .b({_al_u1250_o,_al_u1271_o}),
    .c({_al_u1249_o,_al_u1272_o}),
    .d({_al_u1252_o,_al_u1273_o}),
    .e({_al_u1251_o,\t/a/ID_rs2 [2]}),
    .f({_al_u1253_o,_al_u1274_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1258|t/a/regfile/reg0_b930  (
    .a({_al_u1253_o,_al_u1254_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_4 }),
    .c({_al_u1257_o,\t/a/ID_rs2$1$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1255_o,\t/a/regfile/regfile$28$ [2]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [2]}),
    .mi({open_n1724,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u1258_o,_al_u1255_o}),
    .q({open_n1739,\t/a/regfile/regfile$29$ [2]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100000101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1263|t/a/regfile/reg0_b93  (
    .a({\t/a/ID_rs2$1$_placeOpt_18 ,\t/a/regfile/regfile$2$ [29]}),
    .b({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs1$1$_placeOpt_18 }),
    .c({\t/a/regfile/regfile$3$ [29],\t/a/regfile/regfile$3$ [29]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [29],\t/a/ID_rs1$0$_placeOpt_18 }),
    .mi({open_n1750,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1263_o,_al_u557_o}),
    .q({open_n1754,\t/a/regfile/regfile$2$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1264 (
    .a({_al_u1260_o,_al_u1260_o}),
    .b({_al_u1261_o,_al_u1261_o}),
    .c({_al_u1262_o,_al_u1262_o}),
    .d({_al_u1263_o,_al_u1263_o}),
    .mi({open_n1767,\t/a/ID_rs2$2$_placeOpt_3 }),
    .fx({open_n1772,_al_u1264_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011011100000100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1269|t/a/regfile/reg0_b445  (
    .a({_al_u1266_o,_al_u1265_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_15 }),
    .c({_al_u1268_o,\t/a/ID_rs2$1$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1264_o,\t/a/regfile/regfile$12$ [29]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [29]}),
    .mi({open_n1776,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1269_o,_al_u1266_o}),
    .q({open_n1791,\t/a/regfile/regfile$13$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUT1("(B*~(D*~(1*~(C)*~(A)+1*C*~(A)+~(1)*C*A+1*C*A)))"),
    .INIT_LUT0(16'b1011000000110000),
    .INIT_LUT1(16'b1100010011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1275 (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [2],\t/a/ID_rs2$1$_placeOpt_20 }),
    .c({\t/a/regfile/regfile$31$ [29],\t/a/ID_rs2 [2]}),
    .d({\t/a/ID_rs2$1$_placeOpt_20 ,\t/a/regfile/regfile$31$ [29]}),
    .mi({open_n1804,\t/a/regfile/regfile$30$ [29]}),
    .fx({open_n1809,_al_u1275_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1279|t/a/regfile/reg0_b957  (
    .a({_al_u1276_o,_al_u1275_o}),
    .b({_al_u1274_o,\t/a/ID_rs2$0$_placeOpt_4 }),
    .c({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1278_o,\t/a/regfile/regfile$28$ [29]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [29]}),
    .mi({open_n1813,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1279_o,_al_u1276_o}),
    .q({open_n1828,\t/a/regfile/regfile$29$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+~B*A*C*~D+B*~A*~C*D+B*A*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000110000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1282|t/a/regfile/reg0_b988  (
    .a({open_n1829,\t/a/regfile/regfile$30$ [28]}),
    .b({\t/a/ID_rs2$0$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$31$ [28],\t/a/ID_rs1$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [28],\t/a/regfile/regfile$31$ [28]}),
    .e({\t/a/ID_rs2$1$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_3 }),
    .mi({open_n1831,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1282_o,_al_u580_o}),
    .q({open_n1846,\t/a/regfile/regfile$30$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1000100010001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1290|t/a/regfile/reg0_b700  (
    .a({_al_u1285_o,_al_u1286_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_4 }),
    .c({_al_u1289_o,\t/a/ID_rs2$1$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1287_o,\t/a/regfile/regfile$20$ [28]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [28]}),
    .mi({open_n1848,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1290_o,_al_u1287_o}),
    .q({open_n1863,\t/a/regfile/regfile$21$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*~B*~A*D+~C*~B*A*D"),
    //.LUTG0("~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("C*~B*~A*~D+C*~B*A*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0101000000000000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1291|t/a/regfile/reg0_b188  (
    .a({open_n1864,_al_u1835_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_19 ,open_n1865}),
    .c({\t/a/ID_rs2$0$_placeOpt_19 ,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [28],\t/a/reg_writedat [28]}),
    .e({\t/a/regfile/regfile$4$ [28],\t/a/alu_A_select [1]}),
    .mi({open_n1867,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1291_o,\t/a/aluin/sel0_b28/B0 }),
    .q({open_n1882,\t/a/regfile/regfile$5$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1294|t/a/regfile/reg0_b92  (
    .a({\t/a/ID_rs2$0$_placeOpt_14 ,\t/a/regfile/regfile$2$ [28]}),
    .b({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$3$ [28],\t/a/regfile/regfile$3$ [28]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [28],\t/a/ID_rs1$0$_placeOpt_3 }),
    .mi({open_n1893,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1294_o,_al_u568_o}),
    .q({open_n1897,\t/a/regfile/regfile$2$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1295 (
    .a({_al_u1291_o,_al_u1291_o}),
    .b({_al_u1292_o,_al_u1292_o}),
    .c({_al_u1293_o,_al_u1293_o}),
    .d({_al_u1294_o,_al_u1294_o}),
    .mi({open_n1910,\t/a/ID_rs2$2$_placeOpt_10 }),
    .fx({open_n1915,_al_u1295_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1300|t/a/regfile/reg0_b444  (
    .a({_al_u1295_o,_al_u1296_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_10 }),
    .c({_al_u1299_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1297_o,\t/a/regfile/regfile$12$ [28]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [28]}),
    .mi({open_n1919,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1300_o,_al_u1297_o}),
    .q({open_n1934,\t/a/regfile/regfile$13$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~B*~D*~C*~A+B*~D*~C*~A+~B*D*~C*~A+B*D*~C*~A+~B*~D*C*~A+B*~D*C*~A"),
    //.LUTG0("0"),
    //.LUTG1("~B*~D*C*~A+B*~D*C*~A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0000010101010101),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1302|t/a/regfile/reg0_b187  (
    .a({\t/a/ID_rs2$1$_placeOpt_19 ,open_n1935}),
    .b({open_n1936,\t/a/alu_A_select [1]}),
    .c({\t/a/ID_rs2$0$_placeOpt_19 ,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [27],\t/a/reg_writedat [27]}),
    .e({\t/a/regfile/regfile$4$ [27],_al_u1838_o}),
    .mi({open_n1938,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1302_o,\t/a/aluin/sel0_b27/B0 }),
    .q({open_n1953,\t/a/regfile/regfile$5$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1305|t/a/regfile/reg0_b91  (
    .a({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/regfile/regfile$2$ [27]}),
    .b({\t/a/ID_rs2$1$_placeOpt_12 ,\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/regfile/regfile$3$ [27],\t/a/regfile/regfile$3$ [27]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [27],\t/a/ID_rs1$0$_placeOpt_10 }),
    .mi({open_n1964,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1305_o,_al_u599_o}),
    .q({open_n1968,\t/a/regfile/regfile$2$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1306 (
    .a({_al_u1302_o,_al_u1302_o}),
    .b({_al_u1303_o,_al_u1303_o}),
    .c({_al_u1304_o,_al_u1304_o}),
    .d({_al_u1305_o,_al_u1305_o}),
    .mi({open_n1981,\t/a/ID_rs2$2$_placeOpt_5 }),
    .fx({open_n1986,_al_u1306_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1311|t/a/regfile/reg0_b443  (
    .a({_al_u1306_o,_al_u1307_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_22 }),
    .c({_al_u1310_o,\t/a/ID_rs2$1$_placeOpt_12 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1308_o,\t/a/regfile/regfile$12$ [27]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [27]}),
    .mi({open_n1990,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1311_o,_al_u1308_o}),
    .q({open_n2005,\t/a/regfile/regfile$13$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUT1("(D*~(B*~(1*~(C)*~(A)+1*C*~(A)+~(1)*C*A+1*C*A)))"),
    .INIT_LUT0(16'b1011000000110000),
    .INIT_LUT1(16'b1111011100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1317 (
    .a({\t/a/ID_rs2$0$_placeOpt_16 ,\t/a/ID_rs2$0$_placeOpt_16 }),
    .b({\t/a/ID_rs2$1$_placeOpt_3 ,\t/a/ID_rs2$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$31$ [27],\t/a/ID_rs2$2$_placeOpt_1 }),
    .d({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/regfile/regfile$31$ [27]}),
    .mi({open_n2018,\t/a/regfile/regfile$30$ [27]}),
    .fx({open_n2023,_al_u1317_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1321|t/a/regfile/reg0_b955  (
    .a({_al_u1318_o,_al_u1317_o}),
    .b({_al_u1316_o,\t/a/ID_rs2$0$_placeOpt_16 }),
    .c({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1320_o,\t/a/regfile/regfile$28$ [27]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [27]}),
    .mi({open_n2027,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1321_o,_al_u1318_o}),
    .q({open_n2042,\t/a/regfile/regfile$29$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~C*B*~A*~D+C*B*~A*~D+~C*B*A*~D+C*B*A*~D+C*B*~A*D+C*B*A*D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~C*B*~A*~D+~C*B*A*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b1100000011001100),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1324|t/a/regfile/reg0_b986  (
    .a({open_n2043,\t/a/regfile/regfile$30$ [26]}),
    .b({\t/a/ID_rs2$1$_placeOpt_19 ,\t/a/ID_rs1$1$_placeOpt_15 }),
    .c({\t/a/ID_rs2$0$_placeOpt_19 ,\t/a/ID_rs1$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [26],\t/a/regfile/regfile$31$ [26]}),
    .e({\t/a/regfile/regfile$31$ [26],\t/a/ID_rs1$0$_placeOpt_15 }),
    .mi({open_n2045,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1324_o,_al_u622_o}),
    .q({open_n2060,\t/a/regfile/regfile$30$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100000011000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1332|t/a/regfile/reg0_b698  (
    .a({_al_u1329_o,_al_u1328_o}),
    .b({_al_u1327_o,\t/a/ID_rs2$0$_placeOpt_18 }),
    .c({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1331_o,\t/a/regfile/regfile$20$ [26]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [26]}),
    .mi({open_n2062,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1332_o,_al_u1329_o}),
    .q({open_n2077,\t/a/regfile/regfile$21$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1336|t/a/regfile/reg0_b90  (
    .a({\t/a/ID_rs2$0$_placeOpt_11 ,\t/a/regfile/regfile$2$ [26]}),
    .b({\t/a/ID_rs2$1$_placeOpt_9 ,\t/a/ID_rs1$1$_placeOpt_12 }),
    .c({\t/a/regfile/regfile$3$ [26],\t/a/regfile/regfile$3$ [26]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [26],\t/a/ID_rs1$0$_placeOpt_12 }),
    .mi({open_n2088,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1336_o,_al_u610_o}),
    .q({open_n2092,\t/a/regfile/regfile$2$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1337 (
    .a({_al_u1333_o,_al_u1333_o}),
    .b({_al_u1334_o,_al_u1334_o}),
    .c({_al_u1335_o,_al_u1335_o}),
    .d({_al_u1336_o,_al_u1336_o}),
    .mi({open_n2105,\t/a/ID_rs2$2$_placeOpt_4 }),
    .fx({open_n2110,_al_u1337_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1342|t/a/regfile/reg0_b442  (
    .a({_al_u1337_o,_al_u1338_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_20 }),
    .c({_al_u1341_o,\t/a/ID_rs2$1$_placeOpt_21 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1339_o,\t/a/regfile/regfile$12$ [26]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [26]}),
    .mi({open_n2114,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1342_o,_al_u1339_o}),
    .q({open_n2129,\t/a/regfile/regfile$13$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1347|t/a/regfile/reg0_b89  (
    .a({\t/a/ID_rs2$0$_placeOpt_9 ,\t/a/regfile/regfile$2$ [25]}),
    .b({\t/a/ID_rs2$1$_placeOpt_14 ,\t/a/ID_rs1$1$_placeOpt_21 }),
    .c({\t/a/regfile/regfile$3$ [25],\t/a/regfile/regfile$3$ [25]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [25],\t/a/ID_rs1$0$_placeOpt_21 }),
    .mi({open_n2140,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1347_o,_al_u631_o}),
    .q({open_n2144,\t/a/regfile/regfile$2$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1348 (
    .a({_al_u1344_o,_al_u1344_o}),
    .b({_al_u1345_o,_al_u1345_o}),
    .c({_al_u1346_o,_al_u1346_o}),
    .d({_al_u1347_o,_al_u1347_o}),
    .mi({open_n2157,\t/a/ID_rs2$2$_placeOpt_9 }),
    .fx({open_n2162,_al_u1348_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011011100000100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1353|t/a/regfile/reg0_b441  (
    .a({_al_u1350_o,_al_u1349_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_9 }),
    .c({_al_u1352_o,\t/a/ID_rs2$1$_placeOpt_17 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1348_o,\t/a/regfile/regfile$12$ [25]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [25]}),
    .mi({open_n2166,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1353_o,_al_u1350_o}),
    .q({open_n2181,\t/a/regfile/regfile$13$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1359|t/a/regfile/reg0_b985  (
    .a({\t/a/ID_rs2$0$_placeOpt_19 ,\t/a/regfile/regfile$30$ [25]}),
    .b({\t/a/ID_rs2$1$_placeOpt_14 ,\t/a/ID_rs1$1$_placeOpt_21 }),
    .c({\t/a/ID_rs2$2$_placeOpt_3 ,\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [25],\t/a/regfile/regfile$31$ [25]}),
    .e({\t/a/regfile/regfile$31$ [25],\t/a/ID_rs1$0$_placeOpt_21 }),
    .mi({open_n2183,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1359_o,_al_u643_o}),
    .q({open_n2198,\t/a/regfile/regfile$30$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1363|t/a/regfile/reg0_b953  (
    .a({_al_u1358_o,_al_u1359_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_19 }),
    .c({_al_u1362_o,\t/a/ID_rs2$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1360_o,\t/a/regfile/regfile$28$ [25]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [25]}),
    .mi({open_n2200,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1363_o,_al_u1360_o}),
    .q({open_n2215,\t/a/regfile/regfile$29$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1365|t/a/regfile/reg0_b152  (
    .a({\t/a/ID_rs2$0$_placeOpt_3 ,_al_u2027_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_13 ,\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$4$ [24],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [24],\t/a/reg_writedat [24]}),
    .mi({open_n2226,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1365_o,\t/a/aluin/sel1_b24/B9 }),
    .q({open_n2230,\t/a/regfile/regfile$4$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1368|t/a/regfile/reg0_b88  (
    .a({\t/a/ID_rs2$0$_placeOpt_18 ,\t/a/regfile/regfile$2$ [24]}),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs1$1$_placeOpt_14 }),
    .c({\t/a/regfile/regfile$3$ [24],\t/a/regfile/regfile$3$ [24]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [24],\t/a/ID_rs1$0$_placeOpt_14 }),
    .mi({open_n2241,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1368_o,_al_u652_o}),
    .q({open_n2245,\t/a/regfile/regfile$2$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1374|t/a/regfile/reg0_b440  (
    .a({_al_u1371_o,_al_u1370_o}),
    .b({_al_u1369_o,\t/a/ID_rs2$0$_placeOpt_3 }),
    .c({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_13 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1373_o,\t/a/regfile/regfile$12$ [24]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [24]}),
    .mi({open_n2247,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1374_o,_al_u1371_o}),
    .q({open_n2262,\t/a/regfile/regfile$13$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1379 (
    .a({_al_u1375_o,_al_u1375_o}),
    .b({_al_u1376_o,_al_u1376_o}),
    .c({_al_u1377_o,_al_u1377_o}),
    .d({_al_u1378_o,_al_u1378_o}),
    .mi({open_n2275,\t/a/ID_rs2$2$_placeOpt_9 }),
    .fx({open_n2280,_al_u1379_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1380|t/a/regfile/reg0_b984  (
    .a({\t/a/ID_rs2$0$_placeOpt_19 ,\t/a/regfile/regfile$30$ [24]}),
    .b({\t/a/ID_rs2$1$_placeOpt_14 ,\t/a/ID_rs1$1$_placeOpt_21 }),
    .c({\t/a/ID_rs2$2$_placeOpt_3 ,\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [24],\t/a/regfile/regfile$31$ [24]}),
    .e({\t/a/regfile/regfile$31$ [24],\t/a/ID_rs1$0$_placeOpt_21 }),
    .mi({open_n2284,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1380_o,_al_u664_o}),
    .q({open_n2299,\t/a/regfile/regfile$30$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1384|t/a/regfile/reg0_b952  (
    .a({_al_u1381_o,_al_u1380_o}),
    .b({_al_u1379_o,\t/a/ID_rs2$0$_placeOpt_19 }),
    .c({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_19 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1383_o,\t/a/regfile/regfile$28$ [24]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [24]}),
    .mi({open_n2301,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1384_o,_al_u1381_o}),
    .q({open_n2316,\t/a/regfile/regfile$29$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~C*B*~A*~D+C*B*~A*~D+~C*B*A*~D+C*B*A*~D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~C*B*~A*~D+C*B*~A*~D+~C*B*~A*D+C*B*~A*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0100010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1387|t/a/regfile/reg0_b983  (
    .a({\t/a/regfile/regfile$31$ [23],\t/a/regfile/regfile$30$ [23]}),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({open_n2317,\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [23],\t/a/regfile/regfile$31$ [23]}),
    .e({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .mi({open_n2319,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1387_o,_al_u685_o}),
    .q({open_n2334,\t/a/regfile/regfile$30$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1390|_al_u1579  (
    .a({_al_u1386_o,_al_u1575_o}),
    .b({_al_u1387_o,_al_u1576_o}),
    .c({_al_u1388_o,_al_u1577_o}),
    .d({_al_u1389_o,_al_u1578_o}),
    .e({\t/a/ID_rs2$2$_placeOpt_9 ,\t/a/ID_rs2$2$_placeOpt_9 }),
    .f({_al_u1390_o,_al_u1579_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1000100010001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1395|t/a/regfile/reg0_b695  (
    .a({_al_u1390_o,_al_u1391_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_6 }),
    .c({_al_u1394_o,\t/a/ID_rs2$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1392_o,\t/a/regfile/regfile$20$ [23]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [23]}),
    .mi({open_n2358,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1395_o,_al_u1392_o}),
    .q({open_n2373,\t/a/regfile/regfile$21$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+~A*~B*C*D"),
    //.LUTF1("~A*~C*~D*~B+~A*C*~D*~B+~A*~C*D*~B+~A*C*D*~B+~A*~C*~D*B+~A*~C*D*B"),
    //.LUTG0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("~A*C*~D*~B+~A*C*D*~B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001000000010000),
    .INIT_LUTF1(16'b0001010100010101),
    .INIT_LUTG0(16'b0101000001010000),
    .INIT_LUTG1(16'b0001000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1396|t/a/regfile/reg0_b151  (
    .a({\t/a/ID_rs2$1$_placeOpt_18 ,_al_u2030_o}),
    .b({\t/a/regfile/regfile$5$ [23],\t/a/alu_B_select [1]}),
    .c({\t/a/ID_rs2$0$_placeOpt_15 ,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .e({\t/a/regfile/regfile$4$ [23],\t/a/reg_writedat [23]}),
    .mi({open_n2377,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1396_o,\t/a/aluin/sel1_b23/B9 }),
    .q({open_n2392,\t/a/regfile/regfile$4$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1399|t/a/regfile/reg0_b87  (
    .a({\t/a/ID_rs2$0$_placeOpt_11 ,\t/a/regfile/regfile$2$ [23]}),
    .b({\t/a/ID_rs2$1$_placeOpt_9 ,\t/a/ID_rs1$1$_placeOpt_12 }),
    .c({\t/a/regfile/regfile$3$ [23],\t/a/regfile/regfile$3$ [23]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [23],\t/a/ID_rs1$0$_placeOpt_12 }),
    .mi({open_n2403,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1399_o,_al_u673_o}),
    .q({open_n2407,\t/a/regfile/regfile$2$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1400 (
    .a({_al_u1396_o,_al_u1396_o}),
    .b({_al_u1397_o,_al_u1397_o}),
    .c({_al_u1398_o,_al_u1398_o}),
    .d({_al_u1399_o,_al_u1399_o}),
    .mi({open_n2420,\t/a/ID_rs2$2$_placeOpt_4 }),
    .fx({open_n2425,_al_u1400_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1405|t/a/regfile/reg0_b439  (
    .a({_al_u1400_o,_al_u1401_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_11 }),
    .c({_al_u1404_o,\t/a/ID_rs2$1$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1402_o,\t/a/regfile/regfile$12$ [23]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [23]}),
    .mi({open_n2429,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1405_o,_al_u1402_o}),
    .q({open_n2444,\t/a/regfile/regfile$13$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*~C*~B*D+~A*~C*B*D"),
    //.LUTG0("0"),
    //.LUTG1("A*~C*~B*~D+A*~C*B*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b0000010100001111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1407|t/a/regfile/reg0_b150  (
    .a({\t/a/ID_rs2$0$_placeOpt_3 ,open_n2445}),
    .b({open_n2446,\t/a/alu_B_select [1]}),
    .c({\t/a/ID_rs2$1$_placeOpt_13 ,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [22],\t/a/reg_writedat [22]}),
    .e({\t/a/regfile/regfile$4$ [22],_al_u2033_o}),
    .mi({open_n2448,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1407_o,\t/a/aluin/sel1_b22/B9 }),
    .q({open_n2463,\t/a/regfile/regfile$4$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1410|t/a/regfile/reg0_b86  (
    .a({\t/a/ID_rs2$0$_placeOpt_8 ,\t/a/regfile/regfile$2$ [22]}),
    .b({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$3$ [22],\t/a/regfile/regfile$3$ [22]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [22],\t/a/ID_rs1$0$_placeOpt_3 }),
    .mi({open_n2474,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1410_o,_al_u704_o}),
    .q({open_n2478,\t/a/regfile/regfile$2$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1416|t/a/regfile/reg0_b438  (
    .a({_al_u1413_o,_al_u1412_o}),
    .b({_al_u1411_o,\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1415_o,\t/a/regfile/regfile$12$ [22]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [22]}),
    .mi({open_n2480,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1416_o,_al_u1413_o}),
    .q({open_n2495,\t/a/regfile/regfile$13$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("~D*B*C*~A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1111000011110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1010000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1422|_al_u1674  (
    .a({\t/a/regfile/regfile$31$ [22],\t/a/ID_rs2$0$_placeOpt_14 }),
    .b({\t/a/regfile/regfile$30$ [22],\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/ID_rs2$2$_placeOpt_9 ,\t/a/ID_rs2$2$_placeOpt_9 }),
    .d({\t/a/ID_rs2$0$_placeOpt_14 ,\t/a/regfile/regfile$31$ [11]}),
    .e({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/regfile/regfile$30$ [11]}),
    .f({_al_u1422_o,_al_u1674_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1426|t/a/regfile/reg0_b950  (
    .a({_al_u1421_o,_al_u1422_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_14 }),
    .c({_al_u1425_o,\t/a/ID_rs2$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1423_o,\t/a/regfile/regfile$28$ [22]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [22]}),
    .mi({open_n2519,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1426_o,_al_u1423_o}),
    .q({open_n2534,\t/a/regfile/regfile$29$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+A*B*~C*D+A*B*C*D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*B*~C*~D+~A*B*C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b1000100011001100),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1429|t/a/regfile/reg0_b981  (
    .a({\t/a/ID_rs2$0$_placeOpt_6 ,\t/a/regfile/regfile$30$ [21]}),
    .b({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({open_n2535,\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [21],\t/a/regfile/regfile$31$ [21]}),
    .e({\t/a/regfile/regfile$31$ [21],\t/a/ID_rs1$0$_placeOpt_4 }),
    .mi({open_n2537,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1429_o,_al_u727_o}),
    .q({open_n2552,\t/a/regfile/regfile$30$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1432 (
    .a({_al_u1428_o,_al_u1428_o}),
    .b({_al_u1429_o,_al_u1429_o}),
    .c({_al_u1430_o,_al_u1430_o}),
    .d({_al_u1431_o,_al_u1431_o}),
    .mi({open_n2565,\t/a/ID_rs2$2$_placeOpt_9 }),
    .fx({open_n2570,_al_u1432_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100000011000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1437|t/a/regfile/reg0_b693  (
    .a({_al_u1434_o,_al_u1433_o}),
    .b({_al_u1432_o,\t/a/ID_rs2$0$_placeOpt_6 }),
    .c({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1436_o,\t/a/regfile/regfile$20$ [21]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [21]}),
    .mi({open_n2574,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1437_o,_al_u1434_o}),
    .q({open_n2589,\t/a/regfile/regfile$21$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1438|t/a/regfile/reg0_b149  (
    .a({\t/a/ID_rs2$0$_placeOpt_19 ,_al_u2036_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_19 ,\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$4$ [21],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [21],\t/a/reg_writedat [21]}),
    .mi({open_n2600,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1438_o,\t/a/aluin/sel1_b21/B9 }),
    .q({open_n2604,\t/a/regfile/regfile$4$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1441|t/a/regfile/reg0_b85  (
    .a({\t/a/ID_rs2$0$_placeOpt_17 ,\t/a/regfile/regfile$2$ [21]}),
    .b({\t/a/ID_rs2$1$_placeOpt_8 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$3$ [21],\t/a/regfile/regfile$3$ [21]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [21],\t/a/ID_rs1$0$_placeOpt_11 }),
    .mi({open_n2615,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1441_o,_al_u715_o}),
    .q({open_n2619,\t/a/regfile/regfile$2$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1442 (
    .a({_al_u1438_o,_al_u1438_o}),
    .b({_al_u1439_o,_al_u1439_o}),
    .c({_al_u1440_o,_al_u1440_o}),
    .d({_al_u1441_o,_al_u1441_o}),
    .mi({open_n2632,\t/a/ID_rs2$2$_placeOpt_2 }),
    .fx({open_n2637,_al_u1442_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1447|t/a/regfile/reg0_b437  (
    .a({_al_u1442_o,_al_u1443_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_12 }),
    .c({_al_u1446_o,\t/a/ID_rs2$1$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1444_o,\t/a/regfile/regfile$12$ [21]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [21]}),
    .mi({open_n2641,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1447_o,_al_u1444_o}),
    .q({open_n2656,\t/a/regfile/regfile$13$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*~C*D+~A*B*~C*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000010100000101),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1449|_al_u1453  (
    .a({\t/a/ID_rs2$1$_placeOpt_18 ,_al_u1449_o}),
    .b({open_n2657,_al_u1450_o}),
    .c({\t/a/regfile/regfile$4$ [20],_al_u1451_o}),
    .d({\t/a/regfile/regfile$5$ [20],_al_u1452_o}),
    .e({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs2$2$_placeOpt_3 }),
    .f({_al_u1449_o,_al_u1453_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100000101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1452|t/a/regfile/reg0_b84  (
    .a({\t/a/ID_rs2$1$_placeOpt_9 ,\t/a/regfile/regfile$2$ [20]}),
    .b({\t/a/ID_rs2$0$_placeOpt_11 ,\t/a/ID_rs1$1$_placeOpt_12 }),
    .c({\t/a/regfile/regfile$3$ [20],\t/a/regfile/regfile$3$ [20]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [20],\t/a/ID_rs1$0$_placeOpt_12 }),
    .mi({open_n2690,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1452_o,_al_u746_o}),
    .q({open_n2694,\t/a/regfile/regfile$2$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1458|t/a/regfile/reg0_b436  (
    .a({_al_u1453_o,_al_u1454_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_9 }),
    .c({_al_u1457_o,\t/a/ID_rs2$1$_placeOpt_18 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1455_o,\t/a/regfile/regfile$12$ [20]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [20]}),
    .mi({open_n2696,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1458_o,_al_u1455_o}),
    .q({open_n2711,\t/a/regfile/regfile$13$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1463|_al_u1464  (
    .a({_al_u1459_o,\t/a/ID_rs2$0$_placeOpt_1 }),
    .b({_al_u1460_o,\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({_al_u1461_o,\t/a/ID_rs2$2$_placeOpt_8 }),
    .d({_al_u1462_o,\t/a/regfile/regfile$31$ [20]}),
    .e({\t/a/ID_rs2$2$_placeOpt_8 ,\t/a/regfile/regfile$30$ [20]}),
    .f({_al_u1463_o,_al_u1464_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1468|t/a/regfile/reg0_b948  (
    .a({_al_u1463_o,_al_u1464_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_8 }),
    .c({_al_u1467_o,\t/a/ID_rs2$1$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1465_o,\t/a/regfile/regfile$28$ [20]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [20]}),
    .mi({open_n2735,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1468_o,_al_u1465_o}),
    .q({open_n2750,\t/a/regfile/regfile$29$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~A*~(~0*B)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTG0("~(C*~(D*~A*~(~1*B)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0000001100000011),
    .INIT_LUTG0(16'b0101111100001111),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1470|t/a/regfile/reg0_b161  (
    .a({open_n2751,_al_u2072_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$4$ [1],_al_u2073_o}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [1],\t/a/aluin/n10_lutinv }),
    .e({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/reg_writedat [1]}),
    .mi({open_n2753,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u1470_o,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .q({open_n2768,\t/a/regfile/regfile$5$ [1]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~B*~C)*~((~D*~A))*~(0)+(~B*~C)*(~D*~A)*~(0)+~((~B*~C))*(~D*~A)*0+(~B*~C)*(~D*~A)*0)"),
    //.LUTF1("~B*D*~C*~A+B*D*~C*~A+B*D*C*~A+~B*D*~C*A+B*D*~C*A+B*D*C*A"),
    //.LUTG0("~((~B*~C)*~((~D*~A))*~(1)+(~B*~C)*(~D*~A)*~(1)+~((~B*~C))*(~D*~A)*1+(~B*~C)*(~D*~A)*1)"),
    //.LUTG1("~B*D*~C*~A+~B*D*~C*A"),
    .INIT_LUTF0(16'b1111110011111100),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b1111111110101010),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1471|_al_u1474  (
    .a({open_n2769,_al_u1470_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_21 ,_al_u1473_o}),
    .c({\t/a/regfile/regfile$6$ [1],_al_u1472_o}),
    .d({\t/a/ID_rs2$1$_placeOpt_15 ,_al_u1471_o}),
    .e({\t/a/regfile/regfile$7$ [1],\t/a/ID_rs2$2$_placeOpt_7 }),
    .f({_al_u1471_o,_al_u1474_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000101000111010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1479|t/a/regfile/reg0_b417  (
    .a({_al_u1474_o,_al_u1475_o}),
    .b({_al_u1478_o,\t/a/ID_rs2$0$_placeOpt_21 }),
    .c({\t/a/ID_rs2$3$_placeOpt_3 ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1476_o,\t/a/regfile/regfile$12$ [1]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [1]}),
    .mi({open_n2793,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u1479_o,_al_u1476_o}),
    .q({open_n2808,\t/a/regfile/regfile$13$ [1]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1484 (
    .a({_al_u1480_o,_al_u1480_o}),
    .b({_al_u1481_o,_al_u1481_o}),
    .c({_al_u1482_o,_al_u1482_o}),
    .d({_al_u1483_o,_al_u1483_o}),
    .mi({open_n2821,\t/a/ID_rs2 [2]}),
    .fx({open_n2826,_al_u1484_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1489|t/a/regfile/reg0_b929  (
    .a({_al_u1486_o,_al_u1485_o}),
    .b({_al_u1484_o,\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2$3$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_20 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1488_o,\t/a/regfile/regfile$28$ [1]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [1]}),
    .mi({open_n2830,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u1489_o,_al_u1486_o}),
    .q({open_n2845,\t/a/regfile/regfile$29$ [1]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+D*~B*C*A"),
    //.LUTG0("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("~D*~B*~C*~A+~D*~B*~C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0101010100010001),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1491|t/a/regfile/reg0_b147  (
    .a({open_n2846,_al_u2042_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_19 ,\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$4$ [19],open_n2847}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_19 ,\t/a/reg_writedat [19]}),
    .e({\t/a/regfile/regfile$5$ [19],\t/a/aluin/n10_lutinv }),
    .mi({open_n2849,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1491_o,\t/a/aluin/sel1_b19/B9 }),
    .q({open_n2864,\t/a/regfile/regfile$4$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1494|t/a/regfile/reg0_b83  (
    .a({\t/a/ID_rs2$0$_placeOpt_9 ,\t/a/regfile/regfile$2$ [19]}),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_18 }),
    .c({\t/a/regfile/regfile$3$ [19],\t/a/regfile/regfile$3$ [19]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [19],\t/a/ID_rs1$0$_placeOpt_18 }),
    .mi({open_n2875,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1494_o,_al_u778_o}),
    .q({open_n2879,\t/a/regfile/regfile$2$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1495 (
    .a({_al_u1491_o,_al_u1491_o}),
    .b({_al_u1492_o,_al_u1492_o}),
    .c({_al_u1493_o,_al_u1493_o}),
    .d({_al_u1494_o,_al_u1494_o}),
    .mi({open_n2892,\t/a/ID_rs2$2$_placeOpt_3 }),
    .fx({open_n2897,_al_u1495_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1500|t/a/regfile/reg0_b435  (
    .a({_al_u1495_o,_al_u1496_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_13 }),
    .c({_al_u1499_o,\t/a/ID_rs2$1$_placeOpt_17 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1497_o,\t/a/regfile/regfile$12$ [19]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [19]}),
    .mi({open_n2901,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1500_o,_al_u1497_o}),
    .q({open_n2916,\t/a/regfile/regfile$13$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1506|t/a/regfile/reg0_b979  (
    .a({\t/a/ID_rs2$0$_placeOpt_19 ,\t/a/regfile/regfile$30$ [19]}),
    .b({\t/a/ID_rs2$1$_placeOpt_19 ,\t/a/ID_rs1$1$_placeOpt_15 }),
    .c({\t/a/ID_rs2$2$_placeOpt_6 ,\t/a/ID_rs1$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [19],\t/a/regfile/regfile$31$ [19]}),
    .e({\t/a/regfile/regfile$31$ [19],\t/a/ID_rs1$0$_placeOpt_15 }),
    .mi({open_n2918,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1506_o,_al_u790_o}),
    .q({open_n2933,\t/a/regfile/regfile$30$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1510|t/a/regfile/reg0_b947  (
    .a({_al_u1505_o,_al_u1506_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_14 }),
    .c({_al_u1509_o,\t/a/ID_rs2$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1507_o,\t/a/regfile/regfile$28$ [19]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [19]}),
    .mi({open_n2935,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1510_o,_al_u1507_o}),
    .q({open_n2950,\t/a/regfile/regfile$29$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~D*~B*~A*~C+D*~B*~A*~C+~D*~B*A*~C+D*~B*A*~C+~D*~B*~A*C+~D*~B*A*C"),
    //.LUTG0("~C*~B*~D*~A+~C*~B*D*~A+~C*~B*~D*A+~C*B*~D*A+~C*~B*D*A+~C*B*D*A"),
    //.LUTG1("D*~B*~A*~C+D*~B*A*~C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000101100001011),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1512|t/a/regfile/reg0_b146  (
    .a({open_n2951,\t/a/reg_writedat [18]}),
    .b({\t/a/ID_rs2$1$_placeOpt_19 ,\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$5$ [18],_al_u2045_o}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_19 ,open_n2952}),
    .e({\t/a/regfile/regfile$4$ [18],\t/a/aluin/n10_lutinv }),
    .mi({open_n2954,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1512_o,\t/a/aluin/sel1_b18/B9 }),
    .q({open_n2969,\t/a/regfile/regfile$4$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1515|t/a/regfile/reg0_b82  (
    .a({\t/a/ID_rs2$0$_placeOpt_9 ,\t/a/regfile/regfile$2$ [18]}),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_18 }),
    .c({\t/a/regfile/regfile$3$ [18],\t/a/regfile/regfile$3$ [18]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [18],\t/a/ID_rs1$0$_placeOpt_18 }),
    .mi({open_n2980,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1515_o,_al_u809_o}),
    .q({open_n2984,\t/a/regfile/regfile$2$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011011100000100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1521|t/a/regfile/reg0_b434  (
    .a({_al_u1518_o,_al_u1517_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_9 }),
    .c({_al_u1520_o,\t/a/ID_rs2$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1516_o,\t/a/regfile/regfile$12$ [18]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [18]}),
    .mi({open_n2986,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1521_o,_al_u1518_o}),
    .q({open_n3001,\t/a/regfile/regfile$13$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1526|_al_u1527  (
    .a({_al_u1522_o,\t/a/ID_rs2$0$_placeOpt_7 }),
    .b({_al_u1523_o,\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({_al_u1524_o,\t/a/ID_rs2$2$_placeOpt_8 }),
    .d({_al_u1525_o,\t/a/regfile/regfile$31$ [18]}),
    .e({\t/a/ID_rs2$2$_placeOpt_8 ,\t/a/regfile/regfile$30$ [18]}),
    .f({_al_u1526_o,_al_u1527_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1531|t/a/regfile/reg0_b946  (
    .a({_al_u1526_o,_al_u1527_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_8 }),
    .c({_al_u1530_o,\t/a/ID_rs2$1$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1528_o,\t/a/regfile/regfile$28$ [18]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [18]}),
    .mi({open_n3025,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1531_o,_al_u1528_o}),
    .q({open_n3040,\t/a/regfile/regfile$29$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+A*B*~C*D+A*B*C*D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*B*~C*~D+~A*B*C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b1000100011001100),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1534|t/a/regfile/reg0_b977  (
    .a({\t/a/ID_rs2$0$_placeOpt_19 ,\t/a/regfile/regfile$30$ [17]}),
    .b({\t/a/ID_rs2$1$_placeOpt_19 ,\t/a/ID_rs1$1$_placeOpt_15 }),
    .c({open_n3041,\t/a/ID_rs1$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [17],\t/a/regfile/regfile$31$ [17]}),
    .e({\t/a/regfile/regfile$31$ [17],\t/a/ID_rs1$0$_placeOpt_15 }),
    .mi({open_n3043,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1534_o,_al_u832_o}),
    .q({open_n3058,\t/a/regfile/regfile$30$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1537 (
    .a({_al_u1533_o,_al_u1533_o}),
    .b({_al_u1534_o,_al_u1534_o}),
    .c({_al_u1535_o,_al_u1535_o}),
    .d({_al_u1536_o,_al_u1536_o}),
    .mi({open_n3071,\t/a/ID_rs2$2$_placeOpt_9 }),
    .fx({open_n3076,_al_u1537_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100000011000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1542|t/a/regfile/reg0_b689  (
    .a({_al_u1539_o,_al_u1538_o}),
    .b({_al_u1537_o,\t/a/ID_rs2$0$_placeOpt_18 }),
    .c({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1541_o,\t/a/regfile/regfile$20$ [17]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [17]}),
    .mi({open_n3080,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1542_o,_al_u1539_o}),
    .q({open_n3095,\t/a/regfile/regfile$21$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1543|t/a/regfile/reg0_b945  (
    .a({\t/a/ID_rs2$0$_placeOpt_18 ,\t/a/ID_rs2$0$_placeOpt_18 }),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_5 }),
    .c({\t/a/regfile/regfile$5$ [17],\t/a/regfile/regfile$28$ [17]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$4$ [17],\t/a/regfile/regfile$29$ [17]}),
    .mi({open_n3106,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1543_o,_al_u1533_o}),
    .q({open_n3110,\t/a/regfile/regfile$29$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100000011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1545|t/a/regfile/reg0_b49  (
    .a({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/regfile/regfile$1$ [17]}),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$0$ [17],\t/a/regfile/regfile$0$ [17]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [17],\t/a/ID_rs1$0$_placeOpt_11 }),
    .mi({open_n3121,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1545_o,_al_u819_o}),
    .q({open_n3125,\t/a/regfile/regfile$1$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1546|t/a/regfile/reg0_b81  (
    .a({\t/a/ID_rs2$0$_placeOpt_17 ,\t/a/regfile/regfile$2$ [17]}),
    .b({\t/a/ID_rs2$1$_placeOpt_8 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$3$ [17],\t/a/regfile/regfile$3$ [17]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [17],\t/a/ID_rs1$0$_placeOpt_11 }),
    .mi({open_n3136,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1546_o,_al_u820_o}),
    .q({open_n3140,\t/a/regfile/regfile$2$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1547 (
    .a({_al_u1543_o,_al_u1543_o}),
    .b({_al_u1544_o,_al_u1544_o}),
    .c({_al_u1545_o,_al_u1545_o}),
    .d({_al_u1546_o,_al_u1546_o}),
    .mi({open_n3153,\t/a/ID_rs2$2$_placeOpt_2 }),
    .fx({open_n3158,_al_u1547_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1552|t/a/regfile/reg0_b433  (
    .a({_al_u1549_o,_al_u1548_o}),
    .b({_al_u1547_o,\t/a/ID_rs2$0$_placeOpt_17 }),
    .c({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1551_o,\t/a/regfile/regfile$12$ [17]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [17]}),
    .mi({open_n3162,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1552_o,_al_u1549_o}),
    .q({open_n3177,\t/a/regfile/regfile$13$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1554|t/a/regfile/reg0_b240  (
    .a({\t/a/ID_rs2$0$_placeOpt_9 ,\t/a/ID_rs2$0$_placeOpt_9 }),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs2$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$5$ [16],\t/a/regfile/regfile$6$ [16]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$4$ [16],\t/a/regfile/regfile$7$ [16]}),
    .mi({open_n3188,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1554_o,_al_u1555_o}),
    .q({open_n3192,\t/a/regfile/regfile$7$ [16]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100000011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1556|t/a/regfile/reg0_b48  (
    .a({\t/a/ID_rs2$0$_placeOpt_9 ,\t/a/regfile/regfile$1$ [16]}),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$0$ [16],\t/a/regfile/regfile$0$ [16]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [16],\t/a/ID_rs1$0$_placeOpt_17 }),
    .mi({open_n3203,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1556_o,_al_u850_o}),
    .q({open_n3207,\t/a/regfile/regfile$1$ [16]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1557|t/a/regfile/reg0_b80  (
    .a({\t/a/ID_rs2$0$_placeOpt_13 ,\t/a/regfile/regfile$2$ [16]}),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$3$ [16],\t/a/regfile/regfile$3$ [16]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [16],\t/a/ID_rs1$0$_placeOpt_17 }),
    .mi({open_n3218,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1557_o,_al_u851_o}),
    .q({open_n3222,\t/a/regfile/regfile$2$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011011100000100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1563|t/a/regfile/reg0_b432  (
    .a({_al_u1560_o,_al_u1559_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_20 }),
    .c({_al_u1562_o,\t/a/ID_rs2$1$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1558_o,\t/a/regfile/regfile$12$ [16]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [16]}),
    .mi({open_n3224,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1563_o,_al_u1560_o}),
    .q({open_n3239,\t/a/regfile/regfile$13$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1568|_al_u1610  (
    .a({_al_u1564_o,_al_u1606_o}),
    .b({_al_u1565_o,_al_u1607_o}),
    .c({_al_u1566_o,_al_u1608_o}),
    .d({_al_u1567_o,_al_u1609_o}),
    .e({\t/a/ID_rs2$2$_placeOpt_8 ,\t/a/ID_rs2$2$_placeOpt_8 }),
    .f({_al_u1568_o,_al_u1610_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUT1("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .INIT_LUT0(16'b1011000000110000),
    .INIT_LUT1(16'b1111000001110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1569 (
    .a({\t/a/ID_rs2$0$_placeOpt_8 ,\t/a/ID_rs2$0$_placeOpt_8 }),
    .b({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({\t/a/ID_rs2$2$_placeOpt_8 ,\t/a/ID_rs2$2$_placeOpt_8 }),
    .d({\t/a/regfile/regfile$31$ [16],\t/a/regfile/regfile$31$ [16]}),
    .mi({open_n3274,\t/a/regfile/regfile$30$ [16]}),
    .fx({open_n3279,_al_u1569_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1573|t/a/regfile/reg0_b944  (
    .a({_al_u1570_o,_al_u1569_o}),
    .b({_al_u1568_o,\t/a/ID_rs2$0$_placeOpt_8 }),
    .c({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1572_o,\t/a/regfile/regfile$28$ [16]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [16]}),
    .mi({open_n3283,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1573_o,_al_u1570_o}),
    .q({open_n3298,\t/a/regfile/regfile$29$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~C*B*~A*~D+C*B*~A*~D+~C*B*A*~D+C*B*A*~D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~C*B*~A*~D+C*B*~A*~D+~C*B*~A*D+C*B*~A*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0100010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1576|t/a/regfile/reg0_b975  (
    .a({\t/a/regfile/regfile$31$ [15],\t/a/regfile/regfile$30$ [15]}),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({open_n3299,\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [15],\t/a/regfile/regfile$31$ [15]}),
    .e({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .mi({open_n3301,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1576_o,_al_u874_o}),
    .q({open_n3316,\t/a/regfile/regfile$30$ [15]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1000100010001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1584|t/a/regfile/reg0_b687  (
    .a({_al_u1579_o,_al_u1580_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_19 }),
    .c({_al_u1583_o,\t/a/ID_rs2$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1581_o,\t/a/regfile/regfile$20$ [15]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [15]}),
    .mi({open_n3318,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1584_o,_al_u1581_o}),
    .q({open_n3333,\t/a/regfile/regfile$21$ [15]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100000011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1585|t/a/regfile/reg0_b175  (
    .a({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/regfile/regfile$5$ [15]}),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$4$ [15],\t/a/regfile/regfile$4$ [15]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [15],\t/a/ID_rs1$0$_placeOpt_17 }),
    .mi({open_n3344,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1585_o,_al_u859_o}),
    .q({open_n3348,\t/a/regfile/regfile$5$ [15]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100000011),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1587|t/a/regfile/reg0_b47  (
    .a({\t/a/ID_rs2$1$_placeOpt_21 ,\t/a/regfile/regfile$1$ [15]}),
    .b({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .c({\t/a/regfile/regfile$0$ [15],\t/a/regfile/regfile$0$ [15]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [15],\t/a/ID_rs1$0$_placeOpt_9 }),
    .mi({open_n3359,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1587_o,_al_u861_o}),
    .q({open_n3363,\t/a/regfile/regfile$1$ [15]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1588|t/a/regfile/reg0_b79  (
    .a({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/regfile/regfile$2$ [15]}),
    .b({\t/a/ID_rs2$1$_placeOpt_10 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$3$ [15],\t/a/regfile/regfile$3$ [15]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [15],\t/a/ID_rs1$0$_placeOpt_17 }),
    .mi({open_n3374,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1588_o,_al_u862_o}),
    .q({open_n3378,\t/a/regfile/regfile$2$ [15]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1589 (
    .a({_al_u1585_o,_al_u1585_o}),
    .b({_al_u1586_o,_al_u1586_o}),
    .c({_al_u1587_o,_al_u1587_o}),
    .d({_al_u1588_o,_al_u1588_o}),
    .mi({open_n3391,\t/a/ID_rs2$2$_placeOpt_3 }),
    .fx({open_n3396,_al_u1589_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011011100000100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1594|t/a/regfile/reg0_b431  (
    .a({_al_u1591_o,_al_u1590_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_20 }),
    .c({_al_u1593_o,\t/a/ID_rs2$1$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1589_o,\t/a/regfile/regfile$12$ [15]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [15]}),
    .mi({open_n3400,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1594_o,_al_u1591_o}),
    .q({open_n3415,\t/a/regfile/regfile$13$ [15]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100000011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1596|t/a/regfile/reg0_b174  (
    .a({\t/a/ID_rs2$0$_placeOpt_17 ,\t/a/regfile/regfile$5$ [14]}),
    .b({\t/a/ID_rs2$1$_placeOpt_8 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$4$ [14],\t/a/regfile/regfile$4$ [14]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [14],\t/a/ID_rs1$0$_placeOpt_11 }),
    .mi({open_n3426,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1596_o,_al_u880_o}),
    .q({open_n3430,\t/a/regfile/regfile$5$ [14]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000001100000011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1598|_al_u1516  (
    .a({open_n3431,_al_u1512_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,_al_u1513_o}),
    .c({\t/a/regfile/regfile$0$ [14],_al_u1514_o}),
    .d({\t/a/regfile/regfile$1$ [14],_al_u1515_o}),
    .e({\t/a/ID_rs2$0$_placeOpt_9 ,\t/a/ID_rs2$2$_placeOpt_3 }),
    .f({_al_u1598_o,_al_u1516_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1599|t/a/regfile/reg0_b78  (
    .a({\t/a/ID_rs2$0$_placeOpt_13 ,\t/a/regfile/regfile$2$ [14]}),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$3$ [14],\t/a/regfile/regfile$3$ [14]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [14],\t/a/ID_rs1$0$_placeOpt_17 }),
    .mi({open_n3464,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1599_o,_al_u883_o}),
    .q({open_n3468,\t/a/regfile/regfile$2$ [14]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1600 (
    .a({_al_u1596_o,_al_u1596_o}),
    .b({_al_u1597_o,_al_u1597_o}),
    .c({_al_u1598_o,_al_u1598_o}),
    .d({_al_u1599_o,_al_u1599_o}),
    .mi({open_n3481,\t/a/ID_rs2$2$_placeOpt_3 }),
    .fx({open_n3486,_al_u1600_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011011100000100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1605|t/a/regfile/reg0_b430  (
    .a({_al_u1602_o,_al_u1601_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_17 }),
    .c({_al_u1604_o,\t/a/ID_rs2$1$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1600_o,\t/a/regfile/regfile$12$ [14]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [14]}),
    .mi({open_n3490,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1605_o,_al_u1602_o}),
    .q({open_n3505,\t/a/regfile/regfile$13$ [14]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1611|t/a/regfile/reg0_b974  (
    .a({\t/a/ID_rs2$0$_placeOpt_14 ,\t/a/regfile/regfile$30$ [14]}),
    .b({\t/a/ID_rs2$1$_placeOpt_19 ,\t/a/ID_rs1$1$_placeOpt_15 }),
    .c({\t/a/ID_rs2$2$_placeOpt_6 ,\t/a/ID_rs1$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [14],\t/a/regfile/regfile$31$ [14]}),
    .e({\t/a/regfile/regfile$31$ [14],\t/a/ID_rs1$0$_placeOpt_15 }),
    .mi({open_n3507,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1611_o,_al_u895_o}),
    .q({open_n3522,\t/a/regfile/regfile$30$ [14]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1615|t/a/regfile/reg0_b942  (
    .a({_al_u1610_o,_al_u1611_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_14 }),
    .c({_al_u1614_o,\t/a/ID_rs2$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1612_o,\t/a/regfile/regfile$28$ [14]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [14]}),
    .mi({open_n3524,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1615_o,_al_u1612_o}),
    .q({open_n3539,\t/a/regfile/regfile$29$ [14]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100000011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1617|t/a/regfile/reg0_b173  (
    .a({\t/a/ID_rs2$0$_placeOpt_10 ,\t/a/regfile/regfile$5$ [13]}),
    .b({\t/a/ID_rs2$1$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$4$ [13],\t/a/regfile/regfile$4$ [13]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [13],\t/a/ID_rs1$0$_placeOpt_1 }),
    .mi({open_n3550,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1617_o,_al_u911_o}),
    .q({open_n3554,\t/a/regfile/regfile$5$ [13]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~C*~D)*~((~B*~A))*~(0)+(~C*~D)*(~B*~A)*~(0)+~((~C*~D))*(~B*~A)*0+(~C*~D)*(~B*~A)*0)"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+D*~B*C*A"),
    //.LUTG0("~((~C*~D)*~((~B*~A))*~(1)+(~C*~D)*(~B*~A)*~(1)+~((~C*~D))*(~B*~A)*1+(~C*~D)*(~B*~A)*1)"),
    //.LUTG1("~D*~B*~C*~A+~D*~B*~C*A"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1619|_al_u1621  (
    .a({open_n3555,_al_u1617_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_14 ,_al_u1618_o}),
    .c({\t/a/regfile/regfile$0$ [13],_al_u1620_o}),
    .d({\t/a/ID_rs2$0$_placeOpt_19 ,_al_u1619_o}),
    .e({\t/a/regfile/regfile$1$ [13],\t/a/ID_rs2$2$_placeOpt_3 }),
    .f({_al_u1619_o,_al_u1621_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100000101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1620|t/a/regfile/reg0_b77  (
    .a({\t/a/ID_rs2$1$_placeOpt_18 ,\t/a/regfile/regfile$2$ [13]}),
    .b({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs1$1$_placeOpt_18 }),
    .c({\t/a/regfile/regfile$3$ [13],\t/a/regfile/regfile$3$ [13]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [13],\t/a/ID_rs1$0$_placeOpt_18 }),
    .mi({open_n3588,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1620_o,_al_u914_o}),
    .q({open_n3592,\t/a/regfile/regfile$2$ [13]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011011100000100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1626|t/a/regfile/reg0_b429  (
    .a({_al_u1623_o,_al_u1622_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_9 }),
    .c({_al_u1625_o,\t/a/ID_rs2$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1621_o,\t/a/regfile/regfile$12$ [13]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [13]}),
    .mi({open_n3594,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1626_o,_al_u1623_o}),
    .q({open_n3609,\t/a/regfile/regfile$13$ [13]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1631 (
    .a({_al_u1627_o,_al_u1627_o}),
    .b({_al_u1628_o,_al_u1628_o}),
    .c({_al_u1629_o,_al_u1629_o}),
    .d({_al_u1630_o,_al_u1630_o}),
    .mi({open_n3622,\t/a/ID_rs2$2$_placeOpt_8 }),
    .fx({open_n3627,_al_u1631_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUT1("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .INIT_LUT0(16'b1011000000110000),
    .INIT_LUT1(16'b1111000001110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1632 (
    .a({\t/a/ID_rs2$0$_placeOpt_16 ,\t/a/ID_rs2$0$_placeOpt_16 }),
    .b({\t/a/ID_rs2$1$_placeOpt_16 ,\t/a/ID_rs2$1$_placeOpt_16 }),
    .c({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/ID_rs2$2$_placeOpt_1 }),
    .d({\t/a/regfile/regfile$31$ [13],\t/a/regfile/regfile$31$ [13]}),
    .mi({open_n3642,\t/a/regfile/regfile$30$ [13]}),
    .fx({open_n3647,_al_u1632_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1636|t/a/regfile/reg0_b941  (
    .a({_al_u1633_o,_al_u1632_o}),
    .b({_al_u1631_o,\t/a/ID_rs2$0$_placeOpt_1 }),
    .c({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_16 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1635_o,\t/a/regfile/regfile$28$ [13]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [13]}),
    .mi({open_n3651,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1636_o,_al_u1633_o}),
    .q({open_n3666,\t/a/regfile/regfile$29$ [13]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*~C*D+A*B*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1639|t/a/regfile/reg0_b972  (
    .a({open_n3667,\t/a/regfile/regfile$30$ [12]}),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs1$1$_placeOpt_14 }),
    .c({\t/a/regfile/regfile$31$ [12],\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [12],\t/a/regfile/regfile$31$ [12]}),
    .e({\t/a/ID_rs2$0$_placeOpt_18 ,\t/a/ID_rs1$0$_placeOpt_14 }),
    .mi({open_n3669,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1639_o,_al_u937_o}),
    .q({open_n3684,\t/a/regfile/regfile$30$ [12]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1642 (
    .a({_al_u1638_o,_al_u1638_o}),
    .b({_al_u1639_o,_al_u1639_o}),
    .c({_al_u1640_o,_al_u1640_o}),
    .d({_al_u1641_o,_al_u1641_o}),
    .mi({open_n3697,\t/a/ID_rs2$2$_placeOpt_9 }),
    .fx({open_n3702,_al_u1642_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1000100010001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1647|t/a/regfile/reg0_b684  (
    .a({_al_u1642_o,_al_u1643_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_6 }),
    .c({_al_u1646_o,\t/a/ID_rs2$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1644_o,\t/a/regfile/regfile$20$ [12]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [12]}),
    .mi({open_n3706,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1647_o,_al_u1644_o}),
    .q({open_n3721,\t/a/regfile/regfile$21$ [12]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100000011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1648|t/a/regfile/reg0_b172  (
    .a({\t/a/ID_rs2$0$_placeOpt_13 ,\t/a/regfile/regfile$5$ [12]}),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$4$ [12],\t/a/regfile/regfile$4$ [12]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [12],\t/a/ID_rs1$0$_placeOpt_17 }),
    .mi({open_n3732,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1648_o,_al_u922_o}),
    .q({open_n3736,\t/a/regfile/regfile$5$ [12]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~A)*~((~B*~C))*~(0)+(~D*~A)*(~B*~C)*~(0)+~((~D*~A))*(~B*~C)*0+(~D*~A)*(~B*~C)*0)"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+A*~B*D*~C+~A*~B*~D*C+A*~B*~D*C+A*~B*D*C"),
    //.LUTG0("~((~D*~A)*~((~B*~C))*~(1)+(~D*~A)*(~B*~C)*~(1)+~((~D*~A))*(~B*~C)*1+(~D*~A)*(~B*~C)*1)"),
    //.LUTG1("~A*~B*~D*~C+~A*~B*~D*C"),
    .INIT_LUTF0(16'b1111111110101010),
    .INIT_LUTF1(16'b0010001000110011),
    .INIT_LUTG0(16'b1111110011111100),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1650|_al_u1652  (
    .a({\t/a/ID_rs2$0$_placeOpt_20 ,_al_u1650_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_10 ,_al_u1649_o}),
    .c({open_n3737,_al_u1648_o}),
    .d({\t/a/regfile/regfile$0$ [12],_al_u1651_o}),
    .e({\t/a/regfile/regfile$1$ [12],\t/a/ID_rs2$2$_placeOpt_3 }),
    .f({_al_u1650_o,_al_u1652_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1651|t/a/regfile/reg0_b76  (
    .a({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/regfile/regfile$2$ [12]}),
    .b({\t/a/ID_rs2$1$_placeOpt_10 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .c({\t/a/regfile/regfile$3$ [12],\t/a/regfile/regfile$3$ [12]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [12],\t/a/ID_rs1$0$_placeOpt_9 }),
    .mi({open_n3770,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1651_o,_al_u925_o}),
    .q({open_n3774,\t/a/regfile/regfile$2$ [12]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011011100000100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1657|t/a/regfile/reg0_b428  (
    .a({_al_u1654_o,_al_u1653_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_20 }),
    .c({_al_u1656_o,\t/a/ID_rs2$1$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1652_o,\t/a/regfile/regfile$12$ [12]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [12]}),
    .mi({open_n3776,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1657_o,_al_u1654_o}),
    .q({open_n3791,\t/a/regfile/regfile$13$ [12]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100000011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1659|t/a/regfile/reg0_b171  (
    .a({\t/a/ID_rs2$0$_placeOpt_18 ,\t/a/regfile/regfile$5$ [11]}),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs1$1$_placeOpt_14 }),
    .c({\t/a/regfile/regfile$4$ [11],\t/a/regfile/regfile$4$ [11]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [11],\t/a/ID_rs1$0$_placeOpt_14 }),
    .mi({open_n3802,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u1659_o,_al_u953_o}),
    .q({open_n3806,\t/a/regfile/regfile$5$ [11]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~A)*~((~B*~C))*~(0)+(~D*~A)*(~B*~C)*~(0)+~((~D*~A))*(~B*~C)*0+(~D*~A)*(~B*~C)*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTG0("~((~D*~A)*~((~B*~C))*~(1)+(~D*~A)*(~B*~C)*~(1)+~((~D*~A))*(~B*~C)*1+(~D*~A)*(~B*~C)*1)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    .INIT_LUTF0(16'b1111111110101010),
    .INIT_LUTF1(16'b0000001100000011),
    .INIT_LUTG0(16'b1111110011111100),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1661|_al_u1663  (
    .a({open_n3807,_al_u1661_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,_al_u1660_o}),
    .c({\t/a/regfile/regfile$0$ [11],_al_u1659_o}),
    .d({\t/a/regfile/regfile$1$ [11],_al_u1662_o}),
    .e({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs2$2$_placeOpt_2 }),
    .f({_al_u1661_o,_al_u1663_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1662|t/a/regfile/reg0_b75  (
    .a({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/regfile/regfile$2$ [11]}),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$3$ [11],\t/a/regfile/regfile$3$ [11]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [11],\t/a/ID_rs1$0$_placeOpt_11 }),
    .mi({open_n3840,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u1662_o,_al_u956_o}),
    .q({open_n3844,\t/a/regfile/regfile$2$ [11]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(D*~((~C*~A))*~(B)+D*(~C*~A)*~(B)+~(D)*(~C*~A)*B+D*(~C*~A)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011011100000100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1668|t/a/regfile/reg0_b427  (
    .a({_al_u1665_o,_al_u1664_o}),
    .b({\t/a/ID_rs2 [3],\t/a/ID_rs2$0$_placeOpt_9 }),
    .c({_al_u1667_o,\t/a/ID_rs2$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1663_o,\t/a/regfile/regfile$12$ [11]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [11]}),
    .mi({open_n3846,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u1668_o,_al_u1665_o}),
    .q({open_n3861,\t/a/regfile/regfile$13$ [11]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1673 (
    .a({_al_u1669_o,_al_u1669_o}),
    .b({_al_u1670_o,_al_u1670_o}),
    .c({_al_u1671_o,_al_u1671_o}),
    .d({_al_u1672_o,_al_u1672_o}),
    .mi({open_n3874,\t/a/ID_rs2$2$_placeOpt_8 }),
    .fx({open_n3879,_al_u1673_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1678|t/a/regfile/reg0_b939  (
    .a({_al_u1673_o,_al_u1674_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_14 }),
    .c({_al_u1677_o,\t/a/ID_rs2$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1675_o,\t/a/regfile/regfile$28$ [11]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [11]}),
    .mi({open_n3883,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u1678_o,_al_u1675_o}),
    .q({open_n3898,\t/a/regfile/regfile$29$ [11]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*~C*D+A*B*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b0000110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1681|t/a/regfile/reg0_b970  (
    .a({open_n3899,\t/a/regfile/regfile$30$ [10]}),
    .b({\t/a/ID_rs2$1$_placeOpt_16 ,\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [10],\t/a/ID_rs1$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [10],\t/a/regfile/regfile$31$ [10]}),
    .e({\t/a/ID_rs2$0$_placeOpt_1 ,\t/a/ID_rs1 [0]}),
    .mi({open_n3901,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1681_o,_al_u979_o}),
    .q({open_n3916,\t/a/regfile/regfile$30$ [10]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1684 (
    .a({_al_u1680_o,_al_u1680_o}),
    .b({_al_u1681_o,_al_u1681_o}),
    .c({_al_u1682_o,_al_u1682_o}),
    .d({_al_u1683_o,_al_u1683_o}),
    .mi({open_n3929,\t/a/ID_rs2$2$_placeOpt_8 }),
    .fx({open_n3934,_al_u1684_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1000100010001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1689|t/a/regfile/reg0_b682  (
    .a({_al_u1684_o,_al_u1685_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_2 }),
    .c({_al_u1688_o,\t/a/ID_rs2$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1686_o,\t/a/regfile/regfile$20$ [10]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [10]}),
    .mi({open_n3938,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1689_o,_al_u1686_o}),
    .q({open_n3953,\t/a/regfile/regfile$21$ [10]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100000011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1690|t/a/regfile/reg0_b170  (
    .a({\t/a/ID_rs2$0$_placeOpt_16 ,\t/a/regfile/regfile$5$ [10]}),
    .b({\t/a/ID_rs2$1$_placeOpt_16 ,\t/a/ID_rs1$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$4$ [10],\t/a/regfile/regfile$4$ [10]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [10],\t/a/ID_rs1$0$_placeOpt_2 }),
    .mi({open_n3964,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1690_o,_al_u964_o}),
    .q({open_n3968,\t/a/regfile/regfile$5$ [10]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~C*~D)*~((~B*~A))*~(0)+(~C*~D)*(~B*~A)*~(0)+~((~C*~D))*(~B*~A)*0+(~C*~D)*(~B*~A)*0)"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*~C*~B*D+~A*~C*B*D"),
    //.LUTG0("~((~C*~D)*~((~B*~A))*~(1)+(~C*~D)*(~B*~A)*~(1)+~((~C*~D))*(~B*~A)*1+(~C*~D)*(~B*~A)*1)"),
    //.LUTG1("A*~C*~B*~D+A*~C*B*~D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000010100001111),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1692|_al_u1694  (
    .a({\t/a/ID_rs2$0$_placeOpt_8 ,_al_u1690_o}),
    .b({open_n3969,_al_u1691_o}),
    .c({\t/a/ID_rs2$1$_placeOpt_16 ,_al_u1693_o}),
    .d({\t/a/regfile/regfile$1$ [10],_al_u1692_o}),
    .e({\t/a/regfile/regfile$0$ [10],\t/a/ID_rs2$2$_placeOpt_8 }),
    .f({_al_u1692_o,_al_u1694_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110001000100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1693|t/a/regfile/reg0_b74  (
    .a({\t/a/ID_rs2$0$_placeOpt_8 ,\t/a/regfile/regfile$2$ [10]}),
    .b({\t/a/ID_rs2$1$_placeOpt_16 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$3$ [10],\t/a/regfile/regfile$3$ [10]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [10],\t/a/ID_rs1$0$_placeOpt_3 }),
    .mi({open_n4002,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1693_o,_al_u967_o}),
    .q({open_n4006,\t/a/regfile/regfile$2$ [10]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1699|t/a/regfile/reg0_b426  (
    .a({_al_u1696_o,_al_u1695_o}),
    .b({_al_u1694_o,\t/a/ID_rs2$0$_placeOpt_18 }),
    .c({\t/a/ID_rs2$3$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1698_o,\t/a/regfile/regfile$12$ [10]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [10]}),
    .mi({open_n4008,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1699_o,_al_u1696_o}),
    .q({open_n4023,\t/a/regfile/regfile$13$ [10]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*~C*B*A)"),
    //.LUTF1("~B*~C*~A*~D+B*~C*~A*~D+~B*~C*A*~D+B*~C*A*~D+B*~C*~A*D+B*~C*A*D"),
    //.LUTG0("(~1*D*~C*B*A)"),
    //.LUTG1("~B*~C*~A*~D+~B*~C*A*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000110000001111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1701|t/a/regfile/reg0_b160  (
    .a({open_n4024,_al_u254_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs2$1$_placeOpt_11 ,\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$4$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$5$ [0],\t/a/WB_rd [3]}),
    .mi({open_n4026,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1701_o,\t/a/regfile/mux39_b160_sel_is_3_o }),
    .q({open_n4041,\t/a/regfile/regfile$5$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*C*B*A)"),
    //.LUTF1("~C*B*~A*~D+C*B*~A*~D+~C*B*A*~D+C*B*A*~D+~C*B*~A*D+~C*B*A*D"),
    //.LUTG0("(~1*D*C*B*A)"),
    //.LUTG1("C*B*~A*~D+C*B*A*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1702|t/a/regfile/reg0_b224  (
    .a({open_n4042,_al_u254_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$6$ [0],\t/a/WB_rd [3]}),
    .mi({open_n4044,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1702_o,\t/a/regfile/mux39_b224_sel_is_3_o }),
    .q({open_n4059,\t/a/regfile/regfile$7$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*B*A)"),
    //.LUTF1("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D+C*~B*~A*D+C*~B*A*D"),
    //.LUTG0("(~1*~D*~C*B*A)"),
    //.LUTG1("~C*~B*~A*~D+~C*~B*A*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1703|t/a/regfile/reg0_b32  (
    .a({open_n4060,_al_u254_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$0$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$1$ [0],\t/a/WB_rd [3]}),
    .mi({open_n4062,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1703_o,\t/a/regfile/mux39_b32_sel_is_3_o }),
    .q({open_n4077,\t/a/regfile/regfile$1$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*C*~B*A)"),
    //.LUTF1("~C*B*~A*~D+C*B*~A*~D+~C*B*A*~D+C*B*A*~D+~C*B*~A*D+~C*B*A*D"),
    //.LUTG0("(~1*~D*C*~B*A)"),
    //.LUTG1("C*B*~A*~D+C*B*A*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0000110011001100),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1704|t/a/regfile/reg0_b64  (
    .a({open_n4078,_al_u254_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$3$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$2$ [0],\t/a/WB_rd [3]}),
    .mi({open_n4080,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1704_o,\t/a/regfile/mux39_b64_sel_is_3_o }),
    .q({open_n4095,\t/a/regfile/regfile$2$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*B*A)"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(1*D*~C*B*A)"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1707|t/a/regfile/reg0_b416  (
    .a({_al_u1706_o,_al_u254_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$12$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$13$ [0],\t/a/WB_rd [3]}),
    .mi({open_n4097,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1707_o,\t/a/regfile/mux39_b416_sel_is_3_o }),
    .q({open_n4112,\t/a/regfile/regfile$13$ [0]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUT1("(~D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .INIT_LUT0(16'b0000011100000011),
    .INIT_LUT1(16'b0000000011111011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1708 (
    .a({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/regfile/regfile$10$ [0],\t/a/ID_rs2$2$_placeOpt_7 }),
    .d({\t/a/ID_rs2$2$_placeOpt_7 ,\t/a/regfile/regfile$10$ [0]}),
    .mi({open_n4125,\t/a/regfile/regfile$11$ [0]}),
    .fx({open_n4130,_al_u1708_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUT1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .INIT_LUT0(16'b1010001010100000),
    .INIT_LUT1(16'b1010101010101000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1709 (
    .a({_al_u1708_o,_al_u1708_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/ID_rs2$0$_placeOpt_21 }),
    .c({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .d({\t/a/regfile/regfile$8$ [0],\t/a/regfile/regfile$8$ [0]}),
    .mi({open_n4145,\t/a/regfile/regfile$9$ [0]}),
    .fx({open_n4150,_al_u1709_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1710|_al_u1705  (
    .a({_al_u1705_o,_al_u1701_o}),
    .b({_al_u1707_o,_al_u1702_o}),
    .c({_al_u1709_o,_al_u1703_o}),
    .d({\t/a/ID_rs2$3$_placeOpt_3 ,_al_u1704_o}),
    .e({\t/a/ID_rs2 [4],\t/a/ID_rs2$2$_placeOpt_7 }),
    .f({_al_u1710_o,_al_u1705_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*~C*B*A)"),
    //.LUTF1("~C*~A*~B*~D+C*~A*~B*~D+~C*~A*B*~D+C*~A*B*~D+~C*~A*~B*D+~C*~A*B*D"),
    //.LUTG0("(~1*D*~C*B*A)"),
    //.LUTG1("C*~A*~B*~D+C*~A*B*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000010101010101),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1711|t/a/regfile/reg0_b672  (
    .a({\t/a/ID_rs2$1$_placeOpt_12 ,_al_u256_o}),
    .b({open_n4175,\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$20$ [0],\t/a/WB_rd [3]}),
    .mi({open_n4177,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1711_o,\t/a/regfile/mux39_b672_sel_is_3_o }),
    .q({open_n4192,\t/a/regfile/regfile$21$ [0]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1715 (
    .a({_al_u1711_o,_al_u1711_o}),
    .b({_al_u1712_o,_al_u1712_o}),
    .c({_al_u1713_o,_al_u1713_o}),
    .d({_al_u1714_o,_al_u1714_o}),
    .mi({open_n4205,\t/a/ID_rs2$2$_placeOpt_7 }),
    .fx({open_n4210,_al_u1715_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUT1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUT0(16'b0111000000110000),
    .INIT_LUT1(16'b1111000010110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1716 (
    .a({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/ID_rs2$2$_placeOpt_7 ,\t/a/ID_rs2$2$_placeOpt_7 }),
    .d({\t/a/regfile/regfile$30$ [0],\t/a/regfile/regfile$30$ [0]}),
    .mi({open_n4225,\t/a/regfile/regfile$31$ [0]}),
    .fx({open_n4230,_al_u1716_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*~B*A)"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(1*D*~C*~B*A)"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1717|t/a/regfile/reg0_b896  (
    .a({_al_u1716_o,_al_u256_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs2$1$_placeOpt_11 ,\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$28$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$29$ [0],\t/a/WB_rd [3]}),
    .mi({open_n4234,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1717_o,\t/a/regfile/mux39_b896_sel_is_3_o }),
    .q({open_n4249,\t/a/regfile/regfile$28$ [0]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUT1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .INIT_LUT0(16'b1010001010100000),
    .INIT_LUT1(16'b1010101010101000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1719 (
    .a({_al_u1718_o,_al_u1718_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/ID_rs2$0$_placeOpt_22 }),
    .c({\t/a/ID_rs2$1$_placeOpt_12 ,\t/a/ID_rs2$1$_placeOpt_12 }),
    .d({\t/a/regfile/regfile$24$ [0],\t/a/regfile/regfile$24$ [0]}),
    .mi({open_n4262,\t/a/regfile/regfile$25$ [0]}),
    .fx({open_n4267,_al_u1719_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("~A*~D*~B*~C+~A*D*~B*~C+~A*~D*B*~C+A*~D*B*~C+~A*D*B*~C+A*D*B*~C+~A*~D*~B*C+~A*D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("~A*D*~B*~C+~A*D*B*~C+A*D*B*~C+~A*D*~B*C+~A*D*B*C+A*D*B*C"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1101110111011101),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1101110100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1722|_al_u1723  (
    .a({\t/a/MEM_rd [1],_al_u1722_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/MEM_rd [3]}),
    .c({open_n4270,\t/a/MEM_rd [4]}),
    .d({\t/a/ID_rs2$2$_placeOpt_7 ,\t/a/ID_rs2$3$_placeOpt_3 }),
    .e({\t/a/MEM_rd [2],\t/a/ID_rs2 [4]}),
    .f({_al_u1722_o,_al_u1723_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("(A*C)"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("(A*C)"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b1010000010100000),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b1010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1726|_al_u1725  (
    .a({_al_u1725_o,_al_u1724_o}),
    .b({open_n4293,\t/a/MEM_rd [0]}),
    .c({_al_u1723_o,\t/a/MEM_rd [1]}),
    .d({open_n4296,\t/a/ID_rs2$0$_placeOpt_21 }),
    .e({open_n4297,\t/a/ID_rs2$1$_placeOpt_15 }),
    .f({\t/a/risk_jump/n42_lutinv ,_al_u1725_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~B*~C*~D*~A+~B*C*~D*~A+~B*~C*~D*A+B*~C*~D*A+~B*C*~D*A+B*C*~D*A"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~B*~C*~D*~A+~B*C*~D*~A+~B*~C*D*~A+~B*C*D*~A+~B*~C*~D*A+B*~C*~D*A+~B*C*~D*A+B*C*~D*A+~B*~C*D*A+B*~C*D*A+~B*C*D*A+B*C*D*A"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000010111011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1011101110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1730|_al_u348  (
    .a({\t/a/ID_rs1$1$_placeOpt_20 ,_al_u344_o}),
    .b({\t/a/MEM_rd [1],_al_u345_o}),
    .c({open_n4318,_al_u346_o}),
    .d({\t/a/ID_rs1 [3],_al_u347_o}),
    .e({\t/a/MEM_rd [3],\t/a/ID_rs1$2$_placeOpt_9 }),
    .f({_al_u1730_o,_al_u348_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1731|_al_u1728  (
    .a({_al_u1728_o,_al_u1727_o}),
    .b({_al_u1729_o,\t/a/MEM_rd [0]}),
    .c({_al_u1730_o,\t/a/MEM_rd [2]}),
    .d({\t/a/MEM_rd [4],\t/a/ID_rs1$0$_placeOpt_20 }),
    .e({\t/a/ID_rs1 [4],\t/a/ID_rs1$2$_placeOpt_10 }),
    .f({\t/a/risk_jump/n24_lutinv ,_al_u1728_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(~A*~C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0000010000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1732|t/a/mem_wb/reg1_b5  (
    .a({\t/a/MEM_op [6],_al_u251_o}),
    .b({_al_u251_o,_al_u252_o}),
    .c({\t/a/MEM_op [5],\t/a/MEM_op [5]}),
    .ce(\t/a/ex_mem/n0 ),
    .clk(clock_pad),
    .d({_al_u252_o,\t/a/MEM_op [6]}),
    .mi({open_n4373,\t/a/MEM_op [5]}),
    .f({\t/busarbitration/mux5_b0_sel_is_3_o ,memwrite_cs}),
    .q({open_n4378,\t/a/WB_op [5]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*D*C*~B+A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*D*C*B+A*D*C*B"),
    //.LUTG0("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG1("A*~D*~C*~B+A*D*~C*~B+A*D*C*~B+A*~D*~C*B+A*D*~C*B+A*D*C*B"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111111100001111),
    .INIT_LUTG0(16'b0000001110101010),
    .INIT_LUTG1(16'b1010101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1734|_al_u1720  (
    .a({\t/a/ID_rs2$1$_placeOpt_15 ,_al_u1715_o}),
    .b({open_n4379,_al_u1717_o}),
    .c({\t/a/EX_rd [0],_al_u1719_o}),
    .d({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/ID_rs2$3$_placeOpt_3 }),
    .e({\t/a/EX_rd [1],\t/a/ID_rs2 [4]}),
    .f({_al_u1734_o,_al_u1720_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(0@C)*~(D@B))"),
    //.LUT1("(A*~(1@C)*~(B@D))"),
    .INIT_LUT0(16'b0000100000000010),
    .INIT_LUT1(16'b1000000000100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1735 (
    .a({_al_u1734_o,_al_u1734_o}),
    .b({\t/a/ID_rs2$3$_placeOpt_3 ,\t/a/EX_rd [3]}),
    .c({\t/a/EX_rd [4],\t/a/EX_rd [4]}),
    .d({\t/a/EX_rd [3],\t/a/ID_rs2$3$_placeOpt_3 }),
    .mi({open_n4414,\t/a/ID_rs2 [4]}),
    .fx({open_n4419,_al_u1735_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0@C)*~(D*~B))"),
    //.LUT1("(~A*~(1@D)*~(C*~B))"),
    .INIT_LUT0(16'b0000010000000101),
    .INIT_LUT1(16'b0100010100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1737 (
    .a({_al_u1736_o,_al_u1736_o}),
    .b({\t/a/EX_rd [0],\t/a/EX_rd [0]}),
    .c({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/EX_rd [2]}),
    .d({\t/a/EX_rd [2],\t/a/ID_rs2$0$_placeOpt_21 }),
    .mi({open_n4434,\t/a/ID_rs2$2$_placeOpt_7 }),
    .fx({open_n4439,_al_u1737_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~B*~(D*A)))"),
    //.LUT1("(~B*~D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110000011000000),
    .INIT_LUT1(16'b0000000000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1740|t/a/ex_mem/reg2_b4  (
    .a({_al_u1739_o,_al_u1984_o}),
    .b({\t/a/EX_op [4],\t/a/aluin/n10_lutinv }),
    .c({open_n4442,\t/a/EX_fun3 [1]}),
    .clk(clock_pad),
    .d({\t/a/EX_op [3],\t/a/EX_op [4]}),
    .mi({open_n4454,\t/a/EX_op [4]}),
    .sr(rst_pad),
    .f({_al_u1740_o,\t/a/EX_operation [1]}),
    .q({open_n4458,\t/a/MEM_op [4]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*B*A)"),
    //.LUT1("(~D*~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010001000),
    .INIT_LUT1(16'b0000000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1741|t/a/ex_mem/reg2_b6  (
    .a({\t/a/EX_op [5],_al_u1740_o}),
    .b({open_n4459,\t/a/EX_op [5]}),
    .c({_al_u1740_o,open_n4460}),
    .clk(clock_pad),
    .d({\t/a/EX_op [6],\t/a/EX_op [6]}),
    .mi({open_n4472,\t/a/EX_op [6]}),
    .sr(rst_pad),
    .f({\t/a/aluin/n11_lutinv ,\t/a/aluin/n12_lutinv }),
    .q({open_n4476,\t/a/MEM_op [6]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG0("~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG1("~B*~A*C*~D+B*~A*C*~D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    .INIT_LUTF0(16'b1101110111011101),
    .INIT_LUTF1(16'b1111111101010101),
    .INIT_LUTG0(16'b1101110100000000),
    .INIT_LUTG1(16'b1111000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1744|_al_u1729  (
    .a({\t/a/EX_rd [3],\t/a/MEM_rd [0]}),
    .b({open_n4477,\t/a/ID_rs1$0$_placeOpt_20 }),
    .c({\t/a/ID_rs1$1$_placeOpt_20 ,open_n4478}),
    .d({\t/a/ID_rs1 [3],\t/a/ID_rs1 [3]}),
    .e({\t/a/EX_rd [1],\t/a/MEM_rd [3]}),
    .f({_al_u1744_o,_al_u1729_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A)"),
    //.LUT1("(~(A*~C)*~(~B*D))"),
    .INIT_LUT0(16'b0101000001010000),
    .INIT_LUT1(16'b1100010011110101),
    .MODE("LOGIC"))
    \_al_u1745|_al_u1736  (
    .a({\t/a/ID_rs1 [3],\t/a/EX_rd [1]}),
    .b({\t/a/ID_rs1$2$_placeOpt_10 ,open_n4501}),
    .c({\t/a/EX_rd [3],\t/a/ID_rs2$1$_placeOpt_15 }),
    .d({\t/a/EX_rd [2],open_n4504}),
    .f({_al_u1745_o,_al_u1736_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("(C*A*D*~(0@B))"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("(C*A*D*~(1@B))"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1746|_al_u1743  (
    .a({_al_u1744_o,_al_u1742_o}),
    .b({\t/a/EX_rd [4],\t/a/EX_rd [0]}),
    .c({_al_u1745_o,\t/a/EX_rd [1]}),
    .d({_al_u1743_o,\t/a/ID_rs1$0$_placeOpt_20 }),
    .e({\t/a/ID_rs1 [4],\t/a/ID_rs1$1$_placeOpt_20 }),
    .f({\t/a/risk_jump/n11_lutinv ,_al_u1743_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(~A*~((~D*~B))*~(C)+~A*(~D*~B)*~(C)+~(~A)*(~D*~B)*C+~A*(~D*~B)*C))"),
    //.LUT1("(1*~(~A*~((~D*~B))*~(C)+~A*(~D*~B)*~(C)+~(~A)*(~D*~B)*C+~A*(~D*~B)*C))"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1111101011001010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1749 (
    .a({_al_u1733_o,_al_u1733_o}),
    .b({\t/a/risk_jump/n35_lutinv ,\t/a/risk_jump/n35_lutinv }),
    .c({\t/a/aluin/n11_lutinv ,\t/a/aluin/n11_lutinv }),
    .d({\t/a/risk_jump/n11_lutinv ,\t/a/risk_jump/n11_lutinv }),
    .mi({open_n4557,\t/a/condition/n1_lutinv }),
    .fx({open_n4562,\t/a/condition/n0_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*~(D*A)))"),
    //.LUT1("(~B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0011001000110000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"))
    \_al_u1758|_al_u1779  (
    .a({\t/a/condition/n5 [31],\t/a/condition/n5 [12]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [31],\t/a/ID_jump_addr [12]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*~D+C*~B*A*~D+~C*~B*A*D+C*~B*A*D"),
    //.LUTF1("A*~B*~C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    //.LUTG0("~C*~B*A*~D+C*~B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*~B*A*D+C*~B*A*D"),
    //.LUTG1("A*~B*~C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b0010001000100010),
    .INIT_LUTF1(16'b0010001000100010),
    .INIT_LUTG0(16'b0011001100100010),
    .INIT_LUTG1(16'b0011001100100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1759|_al_u1778  (
    .a({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .e({\t/a/condition/n5 [30],\t/a/condition/n5 [13]}),
    .f({\t/a/ID_jump_addr [30],\t/a/ID_jump_addr [13]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*C*~D+B*~A*C*~D+~B*~A*C*D+B*~A*C*D"),
    //.LUTF1("C*~A*~B*~D+C*~A*B*~D+C*~A*~B*D+C*~A*B*D"),
    //.LUTG0("~B*~A*C*~D+B*~A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D"),
    //.LUTG1("C*~A*~B*~D+C*~A*B*~D+~C*~A*~B*D+C*~A*~B*D+~C*~A*B*D+C*~A*B*D"),
    .INIT_LUTF0(16'b0101000001010000),
    .INIT_LUTF1(16'b0101000001010000),
    .INIT_LUTG0(16'b0101010101010000),
    .INIT_LUTG1(16'b0101010101010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1761|_al_u1777  (
    .a({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .e({\t/a/condition/n5 [29],\t/a/condition/n5 [14]}),
    .f({\t/a/ID_jump_addr [29],\t/a/ID_jump_addr [14]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*~(D*A)))"),
    //.LUT1("(~B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0011001000110000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"))
    \_al_u1762|_al_u1776  (
    .a({\t/a/condition/n5 [28],\t/a/condition/n5 [15]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [28],\t/a/ID_jump_addr [15]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*~(D*A)))"),
    //.LUT1("(~B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0011001000110000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"))
    \_al_u1763|_al_u1775  (
    .a({\t/a/condition/n5 [27],\t/a/condition/n5 [16]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [27],\t/a/ID_jump_addr [16]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*C*~A+D*~B*C*~A+~D*~B*C*A+D*~B*C*A"),
    //.LUTF1("~A*B*~D*~C+A*B*~D*~C+~A*B*~D*C+A*B*~D*C"),
    //.LUTG0("~D*~B*C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*~B*C*A+D*~B*C*A"),
    //.LUTG1("A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C"),
    .INIT_LUTF0(16'b0011000000110000),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b0011001000110010),
    .INIT_LUTG1(16'b0000000011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1764|_al_u1774  (
    .a({\t/a/condition/n5 [26],\t/a/condition/sel1/B2 }),
    .b({\t/a/condition/sel0_b12/B1 ,\t/a/condition/n0_lutinv }),
    .c({open_n4673,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/n0_lutinv ,open_n4676}),
    .e({\t/a/condition/sel1/B2 ,\t/a/condition/n5 [17]}),
    .f({\t/a/ID_jump_addr [26],\t/a/ID_jump_addr [17]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*~D+C*~B*A*~D+~C*~B*A*D+C*~B*A*D"),
    //.LUTF1("A*~B*~C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    //.LUTG0("~C*~B*A*~D+C*~B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*~B*A*D+C*~B*A*D"),
    //.LUTG1("A*~B*~C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b0010001000100010),
    .INIT_LUTF1(16'b0010001000100010),
    .INIT_LUTG0(16'b0011001100100010),
    .INIT_LUTG1(16'b0011001100100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1765|_al_u1773  (
    .a({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .e({\t/a/condition/n5 [25],\t/a/condition/n5 [18]}),
    .f({\t/a/ID_jump_addr [25],\t/a/ID_jump_addr [18]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*~(D*A)))"),
    //.LUT1("(~B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0011001000110000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"))
    \_al_u1766|_al_u1772  (
    .a({\t/a/condition/n5 [24],\t/a/condition/n5 [19]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [24],\t/a/ID_jump_addr [19]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*~(D*A)))"),
    //.LUT1("(~B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0011001000110000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"))
    \_al_u1767|_al_u1770  (
    .a({\t/a/condition/n5 [23],\t/a/condition/n5 [20]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [23],\t/a/ID_jump_addr [20]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*C*~A+D*~B*C*~A+~D*~B*C*A+D*~B*C*A"),
    //.LUTF1("C*~B*~D*~A+C*~B*D*~A+C*~B*~D*A+C*~B*D*A"),
    //.LUTG0("~D*~B*C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*~B*C*A+D*~B*C*A"),
    //.LUTG1("C*~B*~D*~A+C*~B*D*~A+~C*~B*~D*A+C*~B*~D*A+~C*~B*D*A+C*~B*D*A"),
    .INIT_LUTF0(16'b0011000000110000),
    .INIT_LUTF1(16'b0011000000110000),
    .INIT_LUTG0(16'b0011001000110010),
    .INIT_LUTG1(16'b0011001000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1768|_al_u1769  (
    .a({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .e(\t/a/condition/n5 [22:21]),
    .f(\t/a/ID_jump_addr [22:21]));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUT1("(~B*~(~(1*C)*~(D*A)))"),
    .INIT_LUT0(16'b0010001000000000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1771 (
    .a({\t/a/condition/n5 [2],\t/a/condition/n5 [2]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/n1_lutinv ,\t/a/condition/n1_lutinv }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .mi({open_n4797,\t/a/ID_rd [2]}),
    .fx({open_n4802,\t/a/ID_jump_addr [2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUT1("(~B*~(~(1*C)*~(D*A)))"),
    .INIT_LUT0(16'b0010001000000000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1780 (
    .a({\t/a/condition/n5 [11],\t/a/condition/n5 [11]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/n1_lutinv ,\t/a/condition/n1_lutinv }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .mi({open_n4817,\t/a/ID_rd [0]}),
    .fx({open_n4822,\t/a/ID_jump_addr [11]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(~(~D*B)*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b1010111100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1783|t/a/id_ex/reg4_b1  (
    .a({\t/a/EX_rs1 [0],\t/a/aluin/sel1_b16/B9 }),
    .b({\t/a/MEM_rd [1],_al_u2007_o}),
    .c({\t/a/MEM_rd [0],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_rs1 [1],\t/a/EX_rs1 [1]}),
    .mi({open_n4836,\t/a/ID_rs1$1$_placeOpt_20 }),
    .sr(rst_pad),
    .f({_al_u1783_o,\t/a/EX_B [16]}),
    .q({open_n4840,\t/a/EX_rs1 [1]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*D*~C*~A+B*D*~C*~A+~B*D*C*~A+B*D*C*~A+~B*D*~C*A+B*D*~C*A+~B*~D*C*A+B*~D*C*A+~B*D*C*A+B*D*C*A"),
    //.LUTF1("(A*~(0@C)*~(B@D))"),
    //.LUTG0("~B*~D*~C*~A+B*~D*~C*~A+~B*D*~C*~A+B*D*~C*~A+~B*~D*C*~A+B*~D*C*~A+~B*D*C*~A+B*D*C*~A+~B*~D*~C*A+B*~D*~C*A+~B*D*~C*A+B*D*~C*A+~B*~D*C*A+B*~D*C*A+~B*D*C*A+B*D*C*A"),
    //.LUTG1("(A*~(1@C)*~(B@D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110100000),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1111111111111111),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1784|t/a/id_ex/reg4_b4  (
    .a({_al_u1783_o,\t/a/EX_rs1 [4]}),
    .b({\t/a/EX_rs1 [2],open_n4841}),
    .c({\t/a/MEM_rd [4],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_rd [2],_al_u2007_o}),
    .e({\t/a/EX_rs1 [4],\t/a/aluin/sel1_b19/B9 }),
    .mi({open_n4844,\t/a/ID_rs1 [4]}),
    .sr(rst_pad),
    .f({_al_u1784_o,\t/a/EX_B [19]}),
    .q({open_n4859,\t/a/EX_rs1 [4]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~A)"),
    //.LUTF1("(A*~C)"),
    //.LUTG0("(B*~A)"),
    //.LUTG1("(A*~C)"),
    .INIT_LUTF0(16'b0100010001000100),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b0100010001000100),
    .INIT_LUTG1(16'b0000101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1785|_al_u1727  (
    .a({\t/a/EX_rs1 [1],\t/a/MEM_rd [1]}),
    .b({open_n4860,\t/a/ID_rs1$1$_placeOpt_20 }),
    .c({\t/a/MEM_rd [1],open_n4861}),
    .f({_al_u1785_o,_al_u1727_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("(~A*~(0@C)*~(D*~B))"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("(~A*~(1@C)*~(D*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111101010101010),
    .INIT_LUTF1(16'b0000010000000101),
    .INIT_LUTG0(16'b1111111111111111),
    .INIT_LUTG1(16'b0100000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1786|t/a/id_ex/reg4_b3  (
    .a({_al_u1785_o,\t/a/aluin/sel1_b18/B9 }),
    .b({\t/a/MEM_rd [0],open_n4888}),
    .c({\t/a/MEM_rd [3],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_rs1 [0],\t/a/EX_rs1 [3]}),
    .e({\t/a/EX_rs1 [3],_al_u2007_o}),
    .mi({open_n4891,\t/a/ID_rs1 [3]}),
    .sr(rst_pad),
    .f({_al_u1786_o,\t/a/EX_B [18]}),
    .q({open_n4906,\t/a/EX_rs1 [3]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(B*A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(B*A)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1787|_al_u1724  (
    .a({_al_u1784_o,open_n4907}),
    .b({_al_u1786_o,open_n4908}),
    .c({open_n4909,\t/a/ID_rs2$2$_placeOpt_7 }),
    .d({open_n4912,\t/a/MEM_rd [2]}),
    .f({\t/a/n9_lutinv ,_al_u1724_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~D)"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"))
    \_al_u1788|_al_u328  (
    .a({\t/a/EX_rs1 [3],\t/a/WB_rd [1]}),
    .b({\t/a/EX_rs1 [4],open_n4935}),
    .c({\t/a/WB_rd [3],open_n4936}),
    .d({\t/a/WB_rd [4],\t/a/ID_rs1$1$_placeOpt_16 }),
    .f({_al_u1788_o,_al_u328_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(0*~C)*~(~D*B))"),
    //.LUT1("(A*~(1*~C)*~(~D*B))"),
    .INIT_LUT0(16'b1010101000100010),
    .INIT_LUT1(16'b1010000000100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1789 (
    .a({_al_u1788_o,_al_u1788_o}),
    .b({\t/a/EX_rs1 [0],\t/a/EX_rs1 [0]}),
    .c({\t/a/EX_rs1 [1],\t/a/EX_rs1 [1]}),
    .d({\t/a/WB_rd [0],\t/a/WB_rd [0]}),
    .mi({open_n4969,\t/a/WB_rd [1]}),
    .fx({open_n4974,_al_u1789_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*D)"),
    //.LUT1("(~(~C*B)*~(~A*D))"),
    .INIT_LUT0(16'b0101010100000000),
    .INIT_LUT1(16'b1010001011110011),
    .MODE("LOGIC"))
    \_al_u1791|_al_u1043  (
    .a({\t/a/WB_rd [1],\t/a/WB_rd [1]}),
    .b({\t/a/EX_rs1 [4],open_n4977}),
    .c({\t/a/WB_rd [4],open_n4978}),
    .d({\t/a/EX_rs1 [1],\t/a/ID_rs2$1$_placeOpt_15 }),
    .f({_al_u1791_o,_al_u1043_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(C*D*~A*~(0@B))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(C*D*~A*~(1@B))"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b0100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1792|_al_u1790  (
    .a({\t/a/n9_lutinv ,_al_u1789_o}),
    .b({\t/a/EX_rs1 [2],\t/a/EX_rs1 [0]}),
    .c({_al_u1791_o,\t/a/EX_rs1 [3]}),
    .d({_al_u1790_o,\t/a/WB_rd [0]}),
    .e({\t/a/WB_rd [2],\t/a/WB_rd [3]}),
    .f({_al_u1792_o,_al_u1790_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*C)"),
    //.LUT1("(~A*~(D*C*B))"),
    .INIT_LUT0(16'b1010000010100000),
    .INIT_LUT1(16'b0001010101010101),
    .MODE("LOGIC"))
    \_al_u1794|_al_u1795  (
    .a({\t/a/regfile/n46 [0],\t/a/n19 }),
    .b({_al_u1793_o,open_n5021}),
    .c({\t/a/WB_op [0],_al_u1792_o}),
    .d({\t/a/WB_op [1],open_n5024}),
    .f({\t/a/n19 ,\t/a/alu_A_select [1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*~A)"),
    //.LUTF1("~A*~C*~D*~B+~A*C*~D*~B+~A*~C*D*~B+~A*C*D*~B+~A*~C*~D*B+~A*C*~D*B+~A*~C*D*B+~A*C*D*B"),
    //.LUTG0("(~1*~D*~C*~B*~A)"),
    //.LUTG1("~A*~C*~D*~B+~A*C*~D*~B+~A*~C*D*~B+~A*C*D*~B+~A*~C*~D*B+~A*C*~D*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0001000101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1797|t/a/mem_wb/reg2_b4  (
    .a({_al_u1796_o,\t/a/MEM_rd [0]}),
    .b({_al_u251_o,\t/a/MEM_rd [1]}),
    .c({open_n5043,\t/a/MEM_rd [2]}),
    .clk(clock_pad),
    .d({\t/a/MEM_op [5],\t/a/MEM_rd [3]}),
    .e({_al_u252_o,\t/a/MEM_rd [4]}),
    .mi({open_n5046,\t/a/MEM_rd [4]}),
    .sr(rst_pad),
    .f({_al_u1797_o,_al_u1796_o}),
    .q({open_n5061,\t/a/WB_rd [4]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTF1("(~C*A)"),
    //.LUTG0("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG1("(~C*A)"),
    .INIT_LUTF0(16'b1010000010100000),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1798|_al_u1733  (
    .a({_al_u1797_o,\t/a/risk_jump/n42_lutinv }),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .e({open_n5068,\t/a/risk_jump/n24_lutinv }),
    .f({_al_u1798_o,_al_u1733_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1800|t/a/regfile/reg0_b105  (
    .a({\t/a/alu_A_select [1],_al_u2606_o_placeOpt_2}),
    .b({\t/a/alu_A_select [0],_al_u2610_o_placeOpt_2}),
    .c({\t/a/MEM_aludat [9],\t/a/MEM_aludat [9]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [9],\t/a/reg_writedat [9]}),
    .mi({open_n5099,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u1800_o,_al_u2716_o}),
    .q({open_n5103,\t/a/regfile/regfile$3$ [9]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTF1("B*~A*C*D+B*A*C*D"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000011111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000010101010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1802|_al_u1806  (
    .a({open_n5104,\t/a/EX_op [5]}),
    .b({_al_u1801_o,open_n5105}),
    .c({\t/a/EX_op [6],open_n5106}),
    .d({\t/a/EX_op [5],_al_u1802_o}),
    .e({\t/a/EX_op [4],_al_u1803_o}),
    .f({_al_u1802_o,_al_u1806_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~A)"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"))
    \_al_u1804|_al_u1114  (
    .a({_al_u1802_o,\t/a/ID_rs2$0$_placeOpt_15 }),
    .b({open_n5129,\t/a/ID_rs2$1$_placeOpt_9 }),
    .c({open_n5130,\t/a/regfile/regfile$6$ [6]}),
    .d({_al_u1803_o,\t/a/regfile/regfile$7$ [6]}),
    .f({\t/a/aluin/n5_lutinv ,_al_u1114_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~A*~(D*~C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1010111110101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1807|t/a/regfile/reg0_b169  (
    .a({\t/a/aluin/sel0_b9/B0 ,_al_u1800_o}),
    .b({open_n5151,\t/a/alu_A_select [1]}),
    .c({_al_u1806_o,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_memstraddr [9],\t/a/reg_writedat [9]}),
    .mi({open_n5162,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [9],\t/a/aluin/sel0_b9/B0 }),
    .q({open_n5166,\t/a/regfile/regfile$5$ [9]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1808|t/a/regfile/reg0_b104  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [8],\t/a/MEM_aludat [8]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [8],\t/a/reg_writedat [8]}),
    .mi({open_n5177,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u1808_o,_al_u2722_o}),
    .q({open_n5181,\t/a/regfile/regfile$3$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*A*C*~D+B*A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTF1("~(~A*~(D*~B))"),
    //.LUTG0("~B*~A*~C*~D+B*~A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG1("~(~A*~(D*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010110100000),
    .INIT_LUTF1(16'b1011101110101010),
    .INIT_LUTG0(16'b1111010111110101),
    .INIT_LUTG1(16'b1011101110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1810|t/a/id_ex/reg7_b8  (
    .a({\t/a/aluin/sel0_b8/B0 ,\t/a/condition/n0_lutinv }),
    .b({_al_u1806_o,open_n5182}),
    .c({open_n5183,\t/a/ID_memstraddr [8]}),
    .clk(clock_pad),
    .d({\t/a/EX_memstraddr [8],\t/memstraddress [8]}),
    .e({open_n5185,_al_u2807_o}),
    .mi({open_n5187,\t/a/ID_memstraddr [8]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [8],_al_u2815_o}),
    .q({open_n5202,\t/a/EX_memstraddr [8]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D"),
    //.LUTF1("~A*~D*~C*~B+~A*D*~C*~B+~A*~D*~C*B+~A*D*~C*B"),
    //.LUTG0("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*~B*D+~A*C*~B*D"),
    //.LUTG1("~A*~D*~C*~B+~A*D*~C*~B+~A*~D*C*~B+~A*D*C*~B"),
    .INIT_LUTF0(16'b0000000001010101),
    .INIT_LUTF1(16'b0000010100000101),
    .INIT_LUTG0(16'b0001000100010001),
    .INIT_LUTG1(16'b0001000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1811|_al_u1817  (
    .a({\t/a/alu_A_select [1],\t/a/alu_A_select [1]}),
    .b({\t/a/MEM_aludat [7],\t/a/MEM_aludat [5]}),
    .c({\t/a/EX_regdat1 [7],open_n5203}),
    .d({open_n5206,\t/a/EX_regdat1 [5]}),
    .e({\t/a/alu_A_select [0],\t/a/alu_A_select [0]}),
    .f({_al_u1811_o,_al_u1817_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010110100000),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1814|t/a/if_id/reg5_b6  (
    .a({\t/a/alu_A_select [1],\t/busarbitration/n3_placeOpt_2 }),
    .b({\t/a/alu_A_select [0],open_n5227}),
    .c({\t/a/EX_regdat1 [6],\t/memstraddress [6]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [6],\t/a/MEM_aludat [6]}),
    .mi({open_n5238,\t/memstraddress [6]}),
    .sr(rst_pad),
    .f({_al_u1814_o,addr[6]}),
    .q({open_n5242,\t/a/ID_memstraddr [6]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUT1("~(~C*~(D*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111100010),
    .INIT_LUT1(16'b1111010111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1819|t/a/id_ex/reg7_b5  (
    .a({_al_u1806_o,_al_u2807_o}),
    .b({open_n5243,\t/a/condition/n0_lutinv }),
    .c({\t/a/aluin/sel0_b5/B0 ,\t/a/ID_memstraddr [5]}),
    .clk(clock_pad),
    .d({\t/a/EX_memstraddr [5],\t/memstraddress [5]}),
    .mi({open_n5255,\t/a/ID_memstraddr [5]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [5],_al_u2822_o}),
    .q({open_n5259,\t/a/EX_memstraddr [5]}));  // flow_line_reg.v(139)
  EG_PHY_PAD #(
    //.LOCATION("P161"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u182 (
    .ipad(clock),
    .di(clock_pad));  // __top.v(4)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A*~(D*~B))"),
    //.LUT1("(~A*~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000101),
    .INIT_LUT1(16'b0000000101010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1820|t/a/ex_mem/reg4_b4  (
    .a({\t/a/alu_A_select [1],_al_u2541_o}),
    .b({\t/a/EX_regdat1 [4],\t/a/alu/n6 [4]}),
    .c({\t/a/alu_A_select [0],_al_u2547_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [4],_al_u2126_o}),
    .sr(rst_pad),
    .f({_al_u1820_o,\t/a/aludat [4]}),
    .q({open_n5293,\t/a/MEM_aludat [4]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1823|t/a/regfile/reg0_b1023  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_1}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/EX_regdat1 [31],\t/a/MEM_aludat [31]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [31],\t/a/reg_writedat [31]}),
    .mi({open_n5304,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1823_o,_al_u2617_o}),
    .q({open_n5308,\t/a/regfile/regfile$31$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1826|t/a/regfile/reg0_b1022  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_1}),
    .c({\t/a/EX_regdat1 [30],\t/a/MEM_aludat [30]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [30],\t/a/reg_writedat [30]}),
    .mi({open_n5319,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1826_o,_al_u2621_o}),
    .q({open_n5323,\t/a/regfile/regfile$31$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~A*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1011101110101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1828|t/a/regfile/reg0_b190  (
    .a({\t/a/aluin/sel0_b30/B0 ,_al_u1826_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({open_n5324,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_memstraddr [30],\t/a/reg_writedat [30]}),
    .mi({open_n5335,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [30],\t/a/aluin/sel0_b30/B0 }),
    .q({open_n5339,\t/a/regfile/regfile$5$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*~A*~C+D*B*~A*~C+~D*B*A*~C+D*B*A*~C+~D*B*~A*C+~D*B*A*C"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D"),
    //.LUTG0("D*B*~A*~C+D*B*A*~C"),
    //.LUTG1("~A*~B*C*~D+~A*~B*C*D"),
    .INIT_LUTF0(16'b0000110011001100),
    .INIT_LUTF1(16'b0001010100010101),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b0001000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1829|_al_u461  (
    .a({\t/a/alu_A_select [1],open_n5340}),
    .b({\t/a/MEM_aludat [3],\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/alu_A_select [0],\t/a/regfile/regfile$7$ [3]}),
    .d({open_n5343,\t/a/ID_rs1$0$_placeOpt_10 }),
    .e({\t/a/EX_regdat1 [3],\t/a/regfile/regfile$6$ [3]}),
    .f({_al_u1829_o,_al_u461_o}));
  EG_PHY_PAD #(
    //.LOCATION("P136"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u183 (
    .ipad(rst),
    .di(rst_pad));  // __top.v(3)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1832|t/a/regfile/reg0_b1021  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_1}),
    .c({\t/a/MEM_aludat [29],\t/a/MEM_aludat [29]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [29],\t/a/reg_writedat [29]}),
    .mi({open_n5391,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1832_o,_al_u2625_o}),
    .q({open_n5395,\t/a/regfile/regfile$31$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~A*~(D*~C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1010111110101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1834|t/a/regfile/reg0_b189  (
    .a({\t/a/aluin/sel0_b29/B0 ,_al_u1832_o}),
    .b({open_n5396,\t/a/alu_A_select [1]}),
    .c({_al_u1806_o,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_memstraddr [29],\t/a/reg_writedat [29]}),
    .mi({open_n5407,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [29],\t/a/aluin/sel0_b29/B0 }),
    .q({open_n5411,\t/a/regfile/regfile$5$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~C*~(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000000111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1835|t/a/regfile/reg0_b1020  (
    .a({\t/a/MEM_aludat [28],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_1}),
    .c({\t/a/alu_A_select [1],\t/a/MEM_aludat [28]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [28],\t/a/reg_writedat [28]}),
    .mi({open_n5422,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1835_o,_al_u2629_o}),
    .q({open_n5426,\t/a/regfile/regfile$31$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~C*~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000100001101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1838|t/a/regfile/reg0_b1019  (
    .a({\t/a/EX_regdat1 [27],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_1}),
    .c({\t/a/alu_A_select [1],\t/a/MEM_aludat [27]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [27],\t/a/reg_writedat [27]}),
    .mi({open_n5437,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1838_o,_al_u2633_o}),
    .q({open_n5441,\t/a/regfile/regfile$31$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1841|t/a/regfile/reg0_b1018  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_1}),
    .c({\t/a/EX_regdat1 [26],\t/a/MEM_aludat [26]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [26],\t/a/reg_writedat [26]}),
    .mi({open_n5452,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1841_o,_al_u2637_o}),
    .q({open_n5456,\t/a/regfile/regfile$31$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~A*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1011101010111010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1843|t/a/regfile/reg0_b186  (
    .a({\t/a/aluin/sel0_b26/B0 ,_al_u1841_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [26],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({open_n5457,\t/a/reg_writedat [26]}),
    .mi({open_n5468,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [26],\t/a/aluin/sel0_b26/B0 }),
    .q({open_n5472,\t/a/regfile/regfile$5$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~C*~(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000000111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1844|t/a/regfile/reg0_b1017  (
    .a({\t/a/MEM_aludat [25],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_1}),
    .c({\t/a/alu_A_select [1],\t/a/MEM_aludat [25]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [25],\t/a/reg_writedat [25]}),
    .mi({open_n5483,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1844_o,_al_u2641_o}),
    .q({open_n5487,\t/a/regfile/regfile$31$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~A*~(C*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1010101011111010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1846|t/a/regfile/reg0_b185  (
    .a({\t/a/aluin/sel0_b25/B0 ,_al_u1844_o}),
    .b({open_n5488,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [25],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1806_o,\t/a/reg_writedat [25]}),
    .mi({open_n5499,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [25],\t/a/aluin/sel0_b25/B0 }),
    .q({open_n5503,\t/a/regfile/regfile$5$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0001000000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1847|t/a/regfile/reg0_b1016  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_3}),
    .b({\t/a/MEM_aludat [24],_al_u2616_o_placeOpt_1}),
    .c({\t/a/alu_A_select [0],\t/a/MEM_aludat [24]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [24],\t/a/reg_writedat [24]}),
    .mi({open_n5514,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1847_o,_al_u2645_o}),
    .q({open_n5518,\t/a/regfile/regfile$31$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~(~A*~(B*~D))"),
    //.LUTG0("~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("~(~A*~(B*~D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010000),
    .INIT_LUTF1(16'b1010101011101110),
    .INIT_LUTG0(16'b0101000000000000),
    .INIT_LUTG1(16'b1010101011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1849|t/a/regfile/reg0_b184  (
    .a({\t/a/aluin/sel0_b24/B0 ,_al_u1847_o}),
    .b({\t/a/EX_memstraddr [24],open_n5519}),
    .c({open_n5520,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1806_o,\t/a/reg_writedat [24]}),
    .e({open_n5521,\t/a/alu_A_select [1]}),
    .mi({open_n5523,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [24],\t/a/aluin/sel0_b24/B0 }),
    .q({open_n5538,\t/a/regfile/regfile$5$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~C*~(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000000111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1850|t/a/regfile/reg0_b1015  (
    .a({\t/a/MEM_aludat [23],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_1}),
    .c({\t/a/alu_A_select [1],\t/a/MEM_aludat [23]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [23],\t/a/reg_writedat [23]}),
    .mi({open_n5549,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1850_o,_al_u2649_o}),
    .q({open_n5553,\t/a/regfile/regfile$31$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*A*~C+D*~B*A*~C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTF1("~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG0("0"),
    //.LUTG1("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100010),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111111101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1852|t/a/regfile/reg0_b183  (
    .a({_al_u1806_o,\t/a/aluin/n5_lutinv }),
    .b({open_n5554,\t/a/alu_A_select [1]}),
    .c({open_n5555,\t/a/reg_writedat [23]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b23/B0 ,open_n5556}),
    .e({\t/a/EX_memstraddr [23],_al_u1850_o}),
    .mi({open_n5558,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [23],\t/a/aluin/sel0_b23/B0 }),
    .q({open_n5573,\t/a/regfile/regfile$5$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1853|t/a/regfile/reg0_b1014  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_3}),
    .c({\t/a/EX_regdat1 [22],\t/a/MEM_aludat [22]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [22],\t/a/reg_writedat [22]}),
    .mi({open_n5584,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1853_o,_al_u2653_o}),
    .q({open_n5588,\t/a/regfile/regfile$31$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1856|t/a/regfile/reg0_b1013  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_1}),
    .c({\t/a/MEM_aludat [21],\t/a/MEM_aludat [21]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [21],\t/a/reg_writedat [21]}),
    .mi({open_n5599,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1856_o,_al_u2657_o}),
    .q({open_n5603,\t/a/regfile/regfile$31$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~C*~(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000000111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1859|t/a/regfile/reg0_b1012  (
    .a({\t/a/MEM_aludat [20],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_1}),
    .c({\t/a/alu_A_select [1],\t/a/MEM_aludat [20]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [20],\t/a/reg_writedat [20]}),
    .mi({open_n5614,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1859_o,_al_u2661_o}),
    .q({open_n5618,\t/a/regfile/regfile$31$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*~D+C*~B*A*~D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("~(~D*~(A*~C))"),
    //.LUTG0("0"),
    //.LUTG1("~(~D*~(A*~C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b1111111100001010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111111100001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1861|t/a/regfile/reg0_b180  (
    .a({\t/a/EX_memstraddr [20],\t/a/aluin/n5_lutinv }),
    .b({open_n5619,\t/a/alu_A_select [1]}),
    .c({_al_u1806_o,open_n5620}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b20/B0 ,\t/a/reg_writedat [20]}),
    .e({open_n5621,_al_u1859_o}),
    .mi({open_n5623,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [20],\t/a/aluin/sel0_b20/B0 }),
    .q({open_n5638,\t/a/regfile/regfile$5$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(~C*~(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b0000010000000111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1862|t/a/id_ex/reg8_b2  (
    .a({\t/a/MEM_aludat [2],_al_u333_o}),
    .b({\t/a/alu_A_select [0],_al_u532_o}),
    .c({\t/a/alu_A_select [1],_al_u542_o}),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [2],\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u1862_o,\t/a/ID_read_dat1 [2]}),
    .q({open_n5655,\t/a/EX_regdat1 [2]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("~(~A*~(D*~C))"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1010111110101010),
    .MODE("LOGIC"))
    \_al_u1864|_al_u1241  (
    .a({\t/a/aluin/sel0_b2/B0 ,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({open_n5656,\t/a/ID_rs2$1$_placeOpt_11 }),
    .c({_al_u1806_o,\t/a/regfile/regfile$0$ [2]}),
    .d({\t/a/EX_memstraddr [2],\t/a/regfile/regfile$1$ [2]}),
    .f({\t/a/EX_A [2],_al_u1241_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1865|t/a/regfile/reg0_b1011  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_3}),
    .c({\t/a/MEM_aludat [19],\t/a/MEM_aludat [19]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [19],\t/a/reg_writedat [19]}),
    .mi({open_n5687,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1865_o,_al_u2665_o}),
    .q({open_n5691,\t/a/regfile/regfile$31$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1868|t/a/regfile/reg0_b1010  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_3}),
    .c({\t/a/MEM_aludat [18],\t/a/MEM_aludat [18]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [18],\t/a/reg_writedat [18]}),
    .mi({open_n5702,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1868_o,_al_u2669_o}),
    .q({open_n5706,\t/a/regfile/regfile$31$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1871|t/a/regfile/reg0_b1009  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_3}),
    .c({\t/a/MEM_aludat [17],\t/a/MEM_aludat [17]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [17],\t/a/reg_writedat [17]}),
    .mi({open_n5717,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1871_o,_al_u2673_o}),
    .q({open_n5721,\t/a/regfile/regfile$31$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(~A*~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b0001000000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1874|t/a/id_ex/reg8_b16  (
    .a({\t/a/alu_A_select [1],_al_u333_o}),
    .b({\t/a/MEM_aludat [16],_al_u847_o}),
    .c({\t/a/alu_A_select [0],_al_u857_o}),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [16],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1874_o,\t/a/ID_read_dat1 [16]}),
    .q({open_n5738,\t/a/EX_regdat1 [16]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(A*~C))"),
    //.LUT1("~(~D*~(B*~C))"),
    .INIT_LUT0(16'b1111111100001010),
    .INIT_LUT1(16'b1111111100001100),
    .MODE("LOGIC"))
    \_al_u1876|_al_u1891  (
    .a({open_n5739,\t/a/EX_memstraddr [11]}),
    .b({\t/a/EX_memstraddr [16],open_n5740}),
    .c({_al_u1806_o,_al_u1806_o}),
    .d({\t/a/aluin/sel0_b16/B0 ,\t/a/aluin/sel0_b11/B0 }),
    .f({\t/a/EX_A [16],\t/a/EX_A [11]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000101000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1877|t/a/regfile/reg0_b655  (
    .a({\t/a/alu_A_select [1],\t/a/ID_rs1$0$_placeOpt_15 }),
    .b({\t/a/alu_A_select [0],\t/a/ID_rs1$1$_placeOpt_15 }),
    .c({\t/a/EX_regdat1 [15],\t/a/regfile/regfile$20$ [15]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [15],\t/a/regfile/regfile$21$ [15]}),
    .mi({open_n5771,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1877_o,_al_u869_o}),
    .q({open_n5775,\t/a/regfile/regfile$20$ [15]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~B*A*~D*~C+B*A*~D*~C+~B*A*D*~C+B*A*D*~C"),
    //.LUTG0("A*~C*~B*~D+A*~C*B*~D"),
    //.LUTG1("~B*~A*~D*~C+B*~A*~D*~C+~B*A*~D*~C+B*A*~D*~C+~B*~A*D*~C+B*~A*D*~C+~B*A*D*~C+B*A*D*~C+~B*~A*~D*C+B*~A*~D*C+~B*A*~D*C+B*A*~D*C+~B*~A*D*C+B*~A*D*C+~B*A*D*C+B*A*D*C"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b0000000000001010),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1879|_al_u1803  (
    .a({\t/a/EX_memstraddr [15],_al_u1801_o}),
    .c({_al_u1806_o,\t/a/EX_op [3]}),
    .d({open_n5780,\t/a/EX_op [6]}),
    .e({\t/a/aluin/sel0_b15/B0 ,\t/a/EX_op [4]}),
    .f({\t/a/EX_A [15],_al_u1803_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1880|t/a/regfile/reg0_b1006  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_3}),
    .c({\t/a/MEM_aludat [14],\t/a/MEM_aludat [14]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [14],\t/a/reg_writedat [14]}),
    .mi({open_n5811,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1880_o,_al_u2693_o}),
    .q({open_n5815,\t/a/regfile/regfile$31$ [14]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~(~A*~(B*~C))"),
    //.LUTG0("~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("~(~A*~(B*~C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010000),
    .INIT_LUTF1(16'b1010111010101110),
    .INIT_LUTG0(16'b0101000000000000),
    .INIT_LUTG1(16'b1010111010101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1882|t/a/regfile/reg0_b142  (
    .a({\t/a/aluin/sel0_b14/B0 ,_al_u1880_o}),
    .b({\t/a/EX_memstraddr [14],open_n5816}),
    .c({_al_u1806_o,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({open_n5817,\t/a/reg_writedat [14]}),
    .e({open_n5818,\t/a/alu_A_select [1]}),
    .mi({open_n5820,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [14],\t/a/aluin/sel0_b14/B0 }),
    .q({open_n5835,\t/a/regfile/regfile$4$ [14]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1883|t/a/regfile/reg0_b1005  (
    .a({\t/a/alu_A_select [1],_al_u2614_o_placeOpt_3}),
    .b({\t/a/alu_A_select [0],_al_u2616_o_placeOpt_3}),
    .c({\t/a/MEM_aludat [13],\t/a/MEM_aludat [13]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [13],\t/a/reg_writedat [13]}),
    .mi({open_n5846,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1883_o,_al_u2697_o}),
    .q({open_n5850,\t/a/regfile/regfile$31$ [13]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*C*~D+~B*A*C*~D+~B*~A*C*D+~B*A*C*D"),
    //.LUTF1("~(~D*~(A*~C))"),
    //.LUTG0("~B*~A*C*D+~B*A*C*D"),
    //.LUTG1("~(~D*~(A*~C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000000110000),
    .INIT_LUTF1(16'b1111111100001010),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b1111111100001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1885|t/a/regfile/reg0_b141  (
    .a({\t/a/EX_memstraddr [13],open_n5851}),
    .b({open_n5852,_al_u1883_o}),
    .c({_al_u1806_o,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b13/B0 ,\t/a/reg_writedat [13]}),
    .e({open_n5853,\t/a/alu_A_select [1]}),
    .mi({open_n5855,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [13],\t/a/aluin/sel0_b13/B0 }),
    .q({open_n5870,\t/a/regfile/regfile$4$ [13]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D*~(~A*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010110000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1886|t/a/regfile/reg0_b140  (
    .a({\t/a/alu_A_select [1],\t/a/reg_writedat [12]}),
    .b({\t/a/alu_A_select [0],\t/a/alu_A_select [1]}),
    .c({\t/a/MEM_aludat [12],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [12],_al_u1886_o}),
    .mi({open_n5881,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1886_o,\t/a/aluin/sel0_b12/B0 }),
    .q({open_n5885,\t/a/regfile/regfile$4$ [12]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D*~(~A*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010110000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1889|t/a/regfile/reg0_b139  (
    .a({\t/a/alu_A_select [1],\t/a/reg_writedat [11]}),
    .b({\t/a/alu_A_select [0],\t/a/alu_A_select [1]}),
    .c({\t/a/MEM_aludat [11],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [11],_al_u1889_o}),
    .mi({open_n5896,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u1889_o,\t/a/aluin/sel0_b11/B0 }),
    .q({open_n5900,\t/a/regfile/regfile$4$ [11]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D"),
    //.LUTF1("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*~B*A*D+C*~B*A*D"),
    //.LUTG0("B*~A*C*~D+B*A*C*~D"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0010001001110111),
    .INIT_LUTG0(16'b0000000011000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1892|t/a/regfile/reg0_b138  (
    .a({\t/a/alu_A_select [0],open_n5901}),
    .b({\t/a/MEM_aludat [10],\t/a/reg_writedat [10]}),
    .c({open_n5902,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [10],_al_u1892_o}),
    .e({\t/a/alu_A_select [1],\t/a/alu_A_select [1]}),
    .mi({open_n5904,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1892_o,\t/a/aluin/sel0_b10/B0 }),
    .q({open_n5919,\t/a/regfile/regfile$4$ [10]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1895|t/a/id_ex/reg8_b1  (
    .a({\t/a/alu_A_select [1],_al_u333_o}),
    .b({\t/a/alu_A_select [0],_al_u763_o}),
    .c({\t/a/MEM_aludat [1],_al_u773_o}),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [1],\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u1895_o,\t/a/ID_read_dat1 [1]}),
    .q({open_n5936,\t/a/EX_regdat1 [1]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*D)"),
    //.LUT1("~(~D*~(C*~B))"),
    .INIT_LUT0(16'b0011001100000000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"))
    \_al_u1897|_al_u2217  (
    .b({_al_u1806_o,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_memstraddr [1],open_n5939}),
    .d({\t/a/aluin/sel0_b1/B0 ,\t/a/alu/n170_lutinv }),
    .f({\t/a/EX_A [1],\t/a/alu/n202_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1898|t/a/regfile/reg0_b992  (
    .a({\t/a/alu_A_select [1],_al_u2606_o_placeOpt_2}),
    .b({\t/a/alu_A_select [0],_al_u2610_o_placeOpt_2}),
    .c({\t/a/MEM_aludat [0],\t/a/MEM_aludat [0]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [0],\t/a/reg_writedat [0]}),
    .mi({open_n5970,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1898_o,_al_u2758_o}),
    .q({open_n5974,\t/a/regfile/regfile$31$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D"),
    //.LUTG0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("A*~C*B*~D+A*C*B*~D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110101010),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b0000000010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1899|t/a/id_ex/reg7_b0  (
    .a({\t/a/reg_writedat [0],\t/a/EX_memstraddr [0]}),
    .b({\t/a/aluin/n5_lutinv ,open_n5975}),
    .clk(clock_pad),
    .d({_al_u1898_o,\t/a/aluin/sel0_b0/B0 }),
    .e({\t/a/alu_A_select [1],_al_u1806_o}),
    .mi({open_n5980,\t/a/ID_memstraddr [0]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b0/B0 ,\t/a/EX_A [0]}),
    .q({open_n5995,\t/a/EX_memstraddr [0]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*D*~A+C*~B*D*~A+~C*B*D*~A+C*B*D*~A+~C*~B*D*A+C*~B*D*A+~C*B*D*A+C*B*D*A"),
    //.LUTF1("(A*C)"),
    //.LUTG0("~C*~B*~D*A+C*~B*~D*A+~C*~B*D*A+C*~B*D*A"),
    //.LUTG1("(A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b1010000010100000),
    .INIT_LUTG0(16'b0010001000100010),
    .INIT_LUTG1(16'b1010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1901|t/a/mem_wb/reg0_b7  (
    .a({i_data[7],i_data[7]}),
    .b({open_n5996,_al_u1908_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,open_n5997}),
    .clk(clock_pad),
    .d({open_n5999,\t/a/MEM_aludat [7]}),
    .e({open_n6000,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .sr(rst_pad),
    .f({\t/a/mux4_b7/B0_0 ,open_n6015}),
    .q({open_n6019,\t/a/reg_writedat [7]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*(D@C))"),
    //.LUTF1("A*~B*~C*~D+A*~B*~C*D"),
    //.LUTG0("(~1*B*A*(D@C))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100010000000),
    .INIT_LUTF1(16'b0000001000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1902|_al_u1027  (
    .a({\t/a/mux4_b7/B0_0 ,memwrite_cs}),
    .b({\t/a/MEM_fun3 [1],\t/a/MEM_regdat2 [13]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .clk(clock_pad),
    .d({open_n6021,\t/a/MEM_fun3 [1]}),
    .e({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [2]}),
    .mi({o_data[13],o_data[13]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({_al_u1902_o,o_data[13]}),
    .q({\trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D"),
    //.LUTG0("~B*~C*D*~A+B*~C*D*~A"),
    //.LUTG1("~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000010100000000),
    .INIT_LUTG1(16'b1111101011111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1903|_al_u1918  (
    .a({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [2]}),
    .c({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [0]}),
    .d({open_n6041,\t/a/MEM_fun3 [1]}),
    .e({\t/a/MEM_fun3 [1],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .f({_al_u1903_o,_al_u1918_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~A*C*~B+D*~A*C*~B+~D*A*~C*B+D*A*~C*B+~D*~A*C*B+D*~A*C*B+~D*A*C*B+D*A*C*B"),
    //.LUTF1("~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("0"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101100011011000),
    .INIT_LUTF1(16'b1100110000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1904|t/a/if_id/reg2_b2  (
    .a({open_n6062,\t/busarbitration/n3_placeOpt_2 }),
    .b({i_data[9],i_data[9]}),
    .c({open_n6063,\t/busarbitration/instruction [9]}),
    .clk(clock_pad),
    .d({\t/busarbitration/mux5_b0_sel_is_3_o ,open_n6065}),
    .e({_al_u1903_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({_al_u1904_o,open_n6080}),
    .q({open_n6084,\t/a/ID_rd [2]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("0"),
    //.LUTG0("0"),
    //.LUTG1("~A*~B*D*~C+A*~B*D*~C+~A*~B*D*C+A*~B*D*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111110000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0011001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1906|t/a/if_id/reg2_b1  (
    .b({_al_u1903_o,\t/busarbitration/n3_placeOpt_2 }),
    .c({open_n6087,\t/busarbitration/instruction [8]}),
    .clk(clock_pad),
    .d({i_data[8],i_data[8]}),
    .e({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({_al_u1906_o,open_n6103}),
    .q({open_n6107,\t/a/ID_rd [1]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("A*B*~C*~D+A*B*C*~D+A*B*~C*D+A*B*C*D"),
    //.LUTG0("~C*~B*~D*A+C*~B*~D*A+~C*B*~D*A+C*B*~D*A"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b0000000010101010),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1908|_al_u1917  (
    .a({\t/a/MEM_fun3 [2],_al_u1916_o}),
    .b({\t/a/MEM_fun3 [1],open_n6108}),
    .d({open_n6113,\t/a/MEM_fun3 [2]}),
    .e({\t/a/MEM_fun3 [0],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .f({_al_u1908_o,_al_u1917_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*A*(~(B)*C*~(D)+B*~(C)*D))"),
    //.LUTF1("~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("(1*A*(~(B)*C*~(D)+B*~(C)*D))"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0101000000000000),
    .INIT_LUTG0(16'b0000100000100000),
    .INIT_LUTG1(16'b0101010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1916|_al_u1935  (
    .a({\t/a/MEM_fun3 [1],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({open_n6134,\t/a/MEM_fun3 [0]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [1]}),
    .clk(clock_pad),
    .d({i_data[15],\t/a/MEM_fun3 [2]}),
    .e({i_data[7],i_data[15]}),
    .mi({i_data[7],i_data[7]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({_al_u1916_o,_al_u1935_o}),
    .q({\trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~D*~C))"),
    //.LUT1("(A*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010101010000),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1940|_al_u2596  (
    .a({i_data[11],_al_u1903_o}),
    .b({_al_u1903_o,open_n6151}),
    .c({open_n6152,i_data[10]}),
    .clk(clock_pad),
    .d({open_n6154,i_data[12]}),
    .mi({i_data[12],i_data[12]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u1940_o,_al_u2596_o}),
    .q({\trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUTG0("~C*~B*~A*D+C*~B*~A*D+~C*~B*A*D+C*~B*A*D"),
    //.LUTG1("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0001101100011011),
    .INIT_LUTG0(16'b0011001100000000),
    .INIT_LUTG1(16'b0001101100011011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1945|t/a/mem_wb/reg0_b3  (
    .a({\t/busarbitration/n3_placeOpt_2 ,\t/a/MEM_aludat [3]}),
    .b({\t/busarbitration/instruction [3],_al_u1908_o}),
    .c({i_data[3],open_n6168}),
    .clk(clock_pad),
    .d({open_n6170,i_data[3]}),
    .e({open_n6171,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .sr(rst_pad),
    .f({\t/instruction$3$_neg_lutinv ,open_n6186}),
    .q({open_n6190,\t/a/reg_writedat [3]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUT1("~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111001001010000),
    .INIT_LUT1(16'b0000010111110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1946|t/a/mem_wb/reg0_b4  (
    .a({\t/busarbitration/instruction [4],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({open_n6191,_al_u1908_o}),
    .c({\t/busarbitration/n3_placeOpt_2 ,\t/a/MEM_aludat [4]}),
    .clk(clock_pad),
    .d({i_data[4],i_data[4]}),
    .sr(rst_pad),
    .f({\t/instruction$4$_neg_lutinv ,open_n6205}),
    .q({open_n6209,\t/a/reg_writedat [4]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(C*~A*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0001000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1947|t/a/if_id/reg6_b4  (
    .a({\t/instruction$3$_neg_lutinv ,open_n6210}),
    .b({_al_u1944_o,\t/a/if_id/n9 }),
    .c({\t/instruction$4$_neg_lutinv ,open_n6211}),
    .clk(clock_pad),
    .d({open_n6213,\t/instruction$4$_neg_lutinv }),
    .sr(rst_pad),
    .f({_al_u1947_o,open_n6226}),
    .q({open_n6230,\t/a/ID_op [4]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*C*~D+B*~A*C*~D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTF1("~((B*C)*~((0*D))*~(A)+(B*C)*(0*D)*~(A)+~((B*C))*(0*D)*A+(B*C)*(0*D)*A)"),
    //.LUTG0("0"),
    //.LUTG1("~((B*C)*~((1*D))*~(A)+(B*C)*(1*D)*~(A)+~((B*C))*(1*D)*A+(B*C)*(1*D)*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111101001010000),
    .INIT_LUTF1(16'b1011111110111111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1948|t/a/if_id/reg6_b1  (
    .a({\t/busarbitration/n3_placeOpt_2 ,\t/busarbitration/n3_placeOpt_2 }),
    .b({\t/busarbitration/instruction [1],open_n6231}),
    .c({\t/busarbitration/instruction [0],\t/busarbitration/instruction [1]}),
    .clk(clock_pad),
    .d({i_data[1],i_data[1]}),
    .e({i_data[0],\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({_al_u1948_o,open_n6247}),
    .q({open_n6251,\t/a/ID_op [1]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~C*~B*~A*D+C*~B*~A*D+~C*~B*A*D+C*~B*A*D"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b1101110111011101),
    .INIT_LUTG0(16'b0011001100000000),
    .INIT_LUTG1(16'b0001000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1949|t/a/mem_wb/reg0_b2  (
    .a({\t/busarbitration/instruction [2],\t/a/MEM_aludat [2]}),
    .b({\t/busarbitration/n3_placeOpt_2 ,_al_u1908_o}),
    .clk(clock_pad),
    .d({open_n6255,i_data[2]}),
    .e({i_data[2],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .sr(rst_pad),
    .f({\t/instruction$2$_neg_lutinv ,open_n6270}),
    .q({open_n6274,\t/a/reg_writedat [2]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(D*~C*~B*A))"),
    //.LUTF1("~A*B*~C*~D+~A*B*C*~D+~A*B*~C*D+~A*B*C*D"),
    //.LUTG0("(1*~(D*~C*~B*A))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b1111110111111111),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1950|_al_u2805  (
    .a({\t/instruction$2$_neg_lutinv ,_al_u2802_o}),
    .b({_al_u1947_o,_al_u1948_o}),
    .c({open_n6275,_al_u1944_o}),
    .d({open_n6278,\t/instruction$4$_neg_lutinv }),
    .e({_al_u1948_o,\t/a/n0_lutinv }),
    .f({_al_u1950_o,\t/a/n2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("A*~B*C*~D+A*B*C*~D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*B*C*~D+A*B*C*~D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010000010100000),
    .INIT_LUTG0(16'b1111110000110000),
    .INIT_LUTG1(16'b1100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1951|_al_u1955  (
    .a({\t/busarbitration/instruction [29],open_n6299}),
    .b({i_data[29],\t/busarbitration/n3_placeOpt_3 }),
    .c({_al_u1950_o,\t/busarbitration/instruction [25]}),
    .clk(clock_pad),
    .d({open_n6301,i_data[25]}),
    .e({\t/busarbitration/n3_placeOpt_3 ,_al_u1950_o}),
    .mi({open_n6303,i_data[25]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({\t/a/IF_skip_addr [9],\t/a/IF_skip_addr [5]}),
    .q({open_n6318,\trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/ctl_this }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTF1("A*C*~B*D+A*C*B*D"),
    //.LUTG0("~(~A*~(B*(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    //.LUTG1("A*~C*~B*~D+A*~C*B*~D+A*~C*~B*D+A*C*~B*D+A*~C*B*D+A*C*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111010101010),
    .INIT_LUTF1(16'b1010000000000000),
    .INIT_LUTG0(16'b1110111011101010),
    .INIT_LUTG1(16'b1010101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1952|_al_u2083  (
    .a({_al_u1950_o,_al_u2078_o}),
    .b({open_n6319,_al_u2080_o}),
    .c({\t/busarbitration/n3_placeOpt_4 ,\t/busarbitration/n3_placeOpt_4 }),
    .clk(clock_pad),
    .d({i_data[28],\t/busarbitration/instruction [28]}),
    .e({\t/busarbitration/instruction [28],i_data[28]}),
    .mi({i_data[28],i_data[28]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .f({\t/a/IF_skip_addr [8],\t/a/IF_skip_addr [28]}),
    .q({\trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTF1("B*C*~A*D+B*C*A*D"),
    //.LUTG0("~(~A*~(B*(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    //.LUTG1("B*~C*~A*~D+B*~C*A*~D+B*~C*~A*D+B*C*~A*D+B*~C*A*D+B*C*A*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111010101010),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1110111011101010),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1953|_al_u2084  (
    .a({open_n6336,_al_u2078_o}),
    .b({_al_u1950_o,_al_u2080_o}),
    .c({\t/busarbitration/n3_placeOpt_4 ,\t/busarbitration/n3_placeOpt_4 }),
    .clk(clock_pad),
    .d({i_data[27],\t/busarbitration/instruction [27]}),
    .e({\t/busarbitration/instruction [27],i_data[27]}),
    .mi({i_data[27],i_data[27]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .f({\t/a/IF_skip_addr [7],\t/a/IF_skip_addr [27]}),
    .q({\trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D"),
    //.LUTG0("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0001101100011011),
    .INIT_LUTG0(16'b1111010111110101),
    .INIT_LUTG1(16'b0001101100011011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1956|_al_u289  (
    .a({\t/busarbitration/n3_placeOpt_2 ,_al_u251_o}),
    .b({\t/busarbitration/instruction [24],open_n6353}),
    .c({i_data[24],\t/a/MEM_op [6]}),
    .clk(clock_pad),
    .e({open_n6357,_al_u252_o}),
    .mi({i_data[24],i_data[24]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .f({_al_u1956_o,\t/busarbitration/n3 }),
    .q({\trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*A*D)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTG0("~(~B*A*D)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110111111111),
    .INIT_LUTF1(16'b0011001100001111),
    .INIT_LUTG0(16'b1101110111111111),
    .INIT_LUTG1(16'b0011001100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1956|_al_u289_placeOpt_1  (
    .a({open_n6373,_al_u252_o}),
    .b({i_data[24],\t/a/MEM_op [6]}),
    .c({\t/busarbitration/instruction [24],open_n6374}),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,_al_u251_o}),
    .mi({i_data[24],i_data[24]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .f({open_n6390,\t/busarbitration/n3_placeOpt_1 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~C*~B*~A+D*~C*~B*~A+~D*C*~B*~A+D*C*~B*~A+~D*~C*B*~A+D*~C*B*~A+~D*C*B*~A+D*C*B*~A+~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+D*C*~B*A+~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D"),
    //.LUTG0("~D*~C*~B*~A+D*~C*~B*~A+~D*C*~B*~A+D*C*~B*~A+~D*~C*B*~A+D*~C*B*~A+~D*C*B*~A+D*C*B*~A+~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0001101100011011),
    .INIT_LUTG0(16'b1101110111011101),
    .INIT_LUTG1(16'b0001101100011011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1956|_al_u289_placeOpt_2  (
    .a({\t/busarbitration/n3 ,_al_u251_o}),
    .b({\t/busarbitration/instruction [24],\t/a/MEM_op [6]}),
    .c({i_data[24],open_n6396}),
    .clk(clock_pad),
    .e({open_n6400,_al_u252_o}),
    .mi({i_data[24],i_data[24]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .f({open_n6413,\t/busarbitration/n3_placeOpt_2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*~A*~C+D*~B*~A*~C+~D*B*~A*~C+D*B*~A*~C+~D*~B*A*~C+D*~B*A*~C+~D*B*A*~C+D*B*A*~C+~D*~B*~A*C+D*~B*~A*C+~D*B*~A*C+D*B*~A*C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG0("~D*~B*~A*~C+D*~B*~A*~C+~D*B*~A*~C+D*B*~A*~C+~D*~B*A*~C+D*~B*A*~C+~D*B*A*~C+D*B*A*~C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0001000110111011),
    .INIT_LUTG0(16'b1010111110101111),
    .INIT_LUTG1(16'b0001000110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1956|_al_u289_placeOpt_3  (
    .a({\t/busarbitration/n3_placeOpt_2 ,\t/a/MEM_op [6]}),
    .b({\t/busarbitration/instruction [24],open_n6419}),
    .c({open_n6420,_al_u251_o}),
    .clk(clock_pad),
    .d({i_data[24],open_n6422}),
    .e({open_n6423,_al_u252_o}),
    .mi({i_data[24],i_data[24]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .f({open_n6436,\t/busarbitration/n3_placeOpt_3 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~D*~B*~C+A*~D*~B*~C+~A*D*~B*~C+A*D*~B*~C+~A*~D*B*~C+A*~D*B*~C+~A*D*B*~C+A*D*B*~C+~A*~D*~B*C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTG0("~A*~D*~B*~C+A*~D*~B*~C+~A*D*~B*~C+A*D*~B*~C+~A*~D*B*~C+A*~D*B*~C+~A*D*B*~C+A*D*B*~C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0011001101010101),
    .INIT_LUTG0(16'b1100111111001111),
    .INIT_LUTG1(16'b0011001101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1956|_al_u289_placeOpt_4  (
    .a({\t/busarbitration/instruction [24],open_n6442}),
    .b({i_data[24],\t/a/MEM_op [6]}),
    .c({open_n6443,_al_u251_o}),
    .clk(clock_pad),
    .d({\t/busarbitration/n3_placeOpt_2 ,open_n6445}),
    .e({open_n6446,_al_u252_o}),
    .mi({i_data[24],i_data[24]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .f({open_n6459,\t/busarbitration/n3_placeOpt_4 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111111111),
    .INIT_LUTF1(16'b0100011101000111),
    .INIT_LUTG0(16'b1111000011111111),
    .INIT_LUTG1(16'b0100011101000111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1956|_al_u289_placeOpt_5  (
    .a({i_data[24],open_n6465}),
    .b({\t/busarbitration/n3_placeOpt_2 ,open_n6466}),
    .c({\t/busarbitration/instruction [24],\t/a/MEM_op [6]}),
    .clk(clock_pad),
    .d({open_n6468,_al_u251_o}),
    .e({open_n6469,_al_u252_o}),
    .mi({i_data[24],i_data[24]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .f({open_n6482,\t/busarbitration/n3_placeOpt_5 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTF1("0"),
    //.LUTG0("0"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1957|t/a/if_id/reg4_b4  (
    .c({_al_u1956_o,_al_u1956_o}),
    .clk(clock_pad),
    .e({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [4],open_n6509}),
    .q({open_n6513,\t/a/ID_rs2 [4]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(~B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0011000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1959|t/a/if_id/reg4_b3  (
    .b({_al_u1958_o,\t/a/if_id/n9 }),
    .c({_al_u1950_o,open_n6516}),
    .clk(clock_pad),
    .d({open_n6518,_al_u1958_o}),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [3],open_n6531}),
    .q({open_n6535,\t/a/ID_rs2 [3]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A)"),
    //.LUT1("(~A*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b0100010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1959|t/a/if_id/reg4_b3_placeOpt_1  (
    .a({_al_u1958_o,\t/a/if_id/n9 }),
    .b({_al_u1950_o,open_n6536}),
    .c({open_n6537,_al_u1958_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n6558,\t/a/ID_rs2$3$_placeOpt_1 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1959|t/a/if_id/reg4_b3_placeOpt_2  (
    .c({_al_u1958_o,_al_u1958_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n6581,\t/a/ID_rs2$3$_placeOpt_2 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1959|t/a/if_id/reg4_b3_placeOpt_3  (
    .a({_al_u1958_o,\t/a/if_id/n9 }),
    .c({_al_u1950_o,_al_u1958_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n6604,\t/a/ID_rs2$3$_placeOpt_3 }));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~D*~C+A*~B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTG0("~A*~B*~D*~C+A*~B*~D*~C+~A*~B*D*~C+A*~B*D*~C"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111110011),
    .INIT_LUTF1(16'b0011001100110011),
    .INIT_LUTG0(16'b0000001100000011),
    .INIT_LUTG1(16'b0000111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1960|_al_u2117  (
    .b({\t/busarbitration/instruction [22],\t/busarbitration/instruction [16]}),
    .c({i_data[22],\t/busarbitration/n3_placeOpt_3 }),
    .clk(clock_pad),
    .e({\t/busarbitration/n3_placeOpt_3 ,i_data[16]}),
    .mi({i_data[16],i_data[16]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u1960_o,_al_u2117_o}),
    .q({\trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A)"),
    //.LUT1("(~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2  (
    .a({open_n6625,\t/a/if_id/n9 }),
    .b({_al_u1960_o,open_n6626}),
    .clk(clock_pad),
    .d({_al_u1950_o,_al_u1960_o}),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [2],open_n6642}),
    .q({open_n6646,\t/a/ID_rs2 [2]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2_placeOpt_1  (
    .a({_al_u1960_o,open_n6647}),
    .b({open_n6648,\t/a/if_id/n9 }),
    .c({_al_u1950_o,open_n6649}),
    .clk(clock_pad),
    .d({open_n6651,_al_u1960_o}),
    .sr(rst_pad),
    .q({open_n6669,\t/a/ID_rs2$2$_placeOpt_1 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2_placeOpt_10  (
    .b({_al_u1950_o,open_n6672}),
    .c({_al_u1960_o,_al_u1960_o}),
    .clk(clock_pad),
    .d({open_n6674,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n6692,\t/a/ID_rs2$2$_placeOpt_10 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2_placeOpt_2  (
    .b({_al_u1950_o,open_n6695}),
    .c({_al_u1960_o,_al_u1960_o}),
    .clk(clock_pad),
    .d({open_n6697,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n6715,\t/a/ID_rs2$2$_placeOpt_2 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A)"),
    //.LUT1("(~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2_placeOpt_3  (
    .a({open_n6716,\t/a/if_id/n9 }),
    .b({_al_u1960_o,open_n6717}),
    .clk(clock_pad),
    .d({_al_u1950_o,_al_u1960_o}),
    .sr(rst_pad),
    .q({open_n6738,\t/a/ID_rs2$2$_placeOpt_3 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0100010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2_placeOpt_4  (
    .a({_al_u1960_o,_al_u1960_o}),
    .b({_al_u1950_o,open_n6739}),
    .clk(clock_pad),
    .d({open_n6743,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n6761,\t/a/ID_rs2$2$_placeOpt_4 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0011000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2_placeOpt_5  (
    .a({open_n6762,\t/a/if_id/n9 }),
    .b({_al_u1960_o,_al_u1960_o}),
    .c({_al_u1950_o,open_n6763}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n6784,\t/a/ID_rs2$2$_placeOpt_5 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2_placeOpt_6  (
    .a({_al_u1960_o,\t/a/if_id/n9 }),
    .b({open_n6785,_al_u1960_o}),
    .c({_al_u1950_o,open_n6786}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n6807,\t/a/ID_rs2$2$_placeOpt_6 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~A*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0100010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2_placeOpt_7  (
    .a({_al_u1960_o,_al_u1960_o}),
    .b({_al_u1950_o,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n6830,\t/a/ID_rs2$2$_placeOpt_7 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0101010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2_placeOpt_8  (
    .a({_al_u1960_o,_al_u1960_o}),
    .b({open_n6831,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .d({_al_u1950_o,open_n6835}),
    .sr(rst_pad),
    .q({open_n6853,\t/a/ID_rs2$2$_placeOpt_8 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2_placeOpt_9  (
    .a({open_n6854,\t/a/if_id/n9 }),
    .b({_al_u1960_o,_al_u1960_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,open_n6858}),
    .sr(rst_pad),
    .q({open_n6876,\t/a/ID_rs2$2$_placeOpt_9 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0  (
    .c({_al_u1962_o,_al_u1962_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [11],open_n6894}),
    .q({open_n6898,\t/a/ID_rs2 [0]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(~D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000000010101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_1  (
    .a({_al_u1950_o,open_n6899}),
    .b({open_n6900,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .d({_al_u1962_o,_al_u1962_o}),
    .sr(rst_pad),
    .q({open_n6921,\t/a/ID_rs2$0$_placeOpt_1 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_10  (
    .c({_al_u1950_o,_al_u1962_o}),
    .clk(clock_pad),
    .d({_al_u1962_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n6944,\t/a/ID_rs2$0$_placeOpt_10 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(~B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0011000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_11  (
    .b({_al_u1962_o,\t/a/if_id/n9 }),
    .c({_al_u1950_o,open_n6947}),
    .clk(clock_pad),
    .d({open_n6949,_al_u1962_o}),
    .sr(rst_pad),
    .q({open_n6967,\t/a/ID_rs2$0$_placeOpt_11 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_12  (
    .a({_al_u1950_o,open_n6968}),
    .b({_al_u1962_o,_al_u1962_o}),
    .clk(clock_pad),
    .d({open_n6972,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n6990,\t/a/ID_rs2$0$_placeOpt_12 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_13  (
    .a({_al_u1962_o,\t/a/if_id/n9 }),
    .c({_al_u1950_o,open_n6993}),
    .clk(clock_pad),
    .d({open_n6995,_al_u1962_o}),
    .sr(rst_pad),
    .q({open_n7013,\t/a/ID_rs2$0$_placeOpt_13 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_14  (
    .a({_al_u1962_o,_al_u1962_o}),
    .c({_al_u1950_o,open_n7016}),
    .clk(clock_pad),
    .d({open_n7018,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7036,\t/a/ID_rs2$0$_placeOpt_14 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_15  (
    .b({_al_u1950_o,_al_u1962_o}),
    .clk(clock_pad),
    .d({_al_u1962_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7059,\t/a/ID_rs2$0$_placeOpt_15 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B)"),
    //.LUT1("(~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000011),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_16  (
    .b({_al_u1962_o,\t/a/if_id/n9 }),
    .c({open_n7062,_al_u1962_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,open_n7064}),
    .sr(rst_pad),
    .q({open_n7082,\t/a/ID_rs2$0$_placeOpt_16 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A)"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_17  (
    .a({open_n7083,\t/a/if_id/n9 }),
    .c({_al_u1962_o,_al_u1962_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,open_n7087}),
    .sr(rst_pad),
    .q({open_n7105,\t/a/ID_rs2$0$_placeOpt_17 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_18  (
    .b({_al_u1962_o,_al_u1962_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7128,\t/a/ID_rs2$0$_placeOpt_18 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0101010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_19  (
    .a({_al_u1962_o,open_n7129}),
    .c({open_n7132,_al_u1962_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7151,\t/a/ID_rs2$0$_placeOpt_19 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_2  (
    .a({_al_u1962_o,open_n7152}),
    .b({open_n7153,\t/a/if_id/n9 }),
    .c({_al_u1950_o,open_n7154}),
    .clk(clock_pad),
    .d({open_n7156,_al_u1962_o}),
    .sr(rst_pad),
    .q({open_n7174,\t/a/ID_rs2$0$_placeOpt_2 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0101010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_20  (
    .a({_al_u1962_o,_al_u1962_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7197,\t/a/ID_rs2$0$_placeOpt_20 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_21  (
    .b({_al_u1950_o,open_n7200}),
    .c({_al_u1962_o,_al_u1962_o}),
    .clk(clock_pad),
    .d({open_n7202,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7220,\t/a/ID_rs2$0$_placeOpt_21 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0011000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_22  (
    .b({_al_u1962_o,_al_u1962_o}),
    .c({_al_u1950_o,open_n7223}),
    .clk(clock_pad),
    .d({open_n7225,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7243,\t/a/ID_rs2$0$_placeOpt_22 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0101010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_3  (
    .a({_al_u1962_o,open_n7244}),
    .c({open_n7247,_al_u1962_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7266,\t/a/ID_rs2$0$_placeOpt_3 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0011000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_4  (
    .b({_al_u1962_o,_al_u1962_o}),
    .c({_al_u1950_o,open_n7269}),
    .clk(clock_pad),
    .d({open_n7271,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7289,\t/a/ID_rs2$0$_placeOpt_4 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_5  (
    .a({_al_u1950_o,open_n7290}),
    .b({_al_u1962_o,_al_u1962_o}),
    .clk(clock_pad),
    .d({open_n7294,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7312,\t/a/ID_rs2$0$_placeOpt_5 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0100010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_6  (
    .a({_al_u1962_o,_al_u1962_o}),
    .b({_al_u1950_o,open_n7313}),
    .clk(clock_pad),
    .d({open_n7317,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7335,\t/a/ID_rs2$0$_placeOpt_6 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B)"),
    //.LUT1("(~C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000011),
    .INIT_LUT1(16'b0000101000001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_7  (
    .a({_al_u1950_o,open_n7336}),
    .b({open_n7337,\t/a/if_id/n9 }),
    .c({_al_u1962_o,_al_u1962_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n7358,\t/a/ID_rs2$0$_placeOpt_7 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_8  (
    .a({_al_u1962_o,_al_u1962_o}),
    .b({open_n7359,\t/a/if_id/n9 }),
    .c({_al_u1950_o,open_n7360}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n7381,\t/a/ID_rs2$0$_placeOpt_8 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(~D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0_placeOpt_9  (
    .b({open_n7384,\t/a/if_id/n9 }),
    .c({_al_u1950_o,open_n7385}),
    .clk(clock_pad),
    .d({_al_u1962_o,_al_u1962_o}),
    .sr(rst_pad),
    .q({open_n7404,\t/a/ID_rs2$0$_placeOpt_9 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1  (
    .b({_al_u1950_o,open_n7407}),
    .c({_al_u1965_o,_al_u1965_o}),
    .clk(clock_pad),
    .d({open_n7409,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [1],open_n7422}),
    .q({open_n7426,\t/a/ID_rs2 [1]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(~D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000000010101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_1  (
    .a({_al_u1950_o,open_n7427}),
    .b({open_n7428,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .d({_al_u1965_o,_al_u1965_o}),
    .sr(rst_pad),
    .q({open_n7449,\t/a/ID_rs2$1$_placeOpt_1 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0101010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_10  (
    .a({_al_u1965_o,_al_u1965_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7472,\t/a/ID_rs2$1$_placeOpt_10 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A)"),
    //.LUT1("(~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_11  (
    .a({_al_u1950_o,\t/a/if_id/n9 }),
    .b({_al_u1965_o,open_n7473}),
    .c({open_n7474,_al_u1965_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n7495,\t/a/ID_rs2$1$_placeOpt_11 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0101010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_12  (
    .a({_al_u1965_o,_al_u1965_o}),
    .b({open_n7496,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .d({_al_u1950_o,open_n7500}),
    .sr(rst_pad),
    .q({open_n7518,\t/a/ID_rs2$1$_placeOpt_12 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_13  (
    .a({_al_u1965_o,_al_u1965_o}),
    .c({_al_u1950_o,open_n7521}),
    .clk(clock_pad),
    .d({open_n7523,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7541,\t/a/ID_rs2$1$_placeOpt_13 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_14  (
    .a({_al_u1950_o,open_n7542}),
    .b({_al_u1965_o,_al_u1965_o}),
    .clk(clock_pad),
    .d({open_n7546,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7564,\t/a/ID_rs2$1$_placeOpt_14 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_15  (
    .c({_al_u1965_o,_al_u1965_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7587,\t/a/ID_rs2$1$_placeOpt_15 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000011),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_16  (
    .a({_al_u1965_o,open_n7588}),
    .b({open_n7589,\t/a/if_id/n9 }),
    .c({_al_u1950_o,_al_u1965_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n7610,\t/a/ID_rs2$1$_placeOpt_16 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_17  (
    .a({_al_u1965_o,\t/a/if_id/n9 }),
    .c({_al_u1950_o,_al_u1965_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n7633,\t/a/ID_rs2$1$_placeOpt_17 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0011000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_18  (
    .b({_al_u1965_o,_al_u1965_o}),
    .c({_al_u1950_o,open_n7636}),
    .clk(clock_pad),
    .d({open_n7638,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7656,\t/a/ID_rs2$1$_placeOpt_18 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_19  (
    .a({_al_u1965_o,_al_u1965_o}),
    .c({_al_u1950_o,open_n7659}),
    .clk(clock_pad),
    .d({open_n7661,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7679,\t/a/ID_rs2$1$_placeOpt_19 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_2  (
    .a({_al_u1950_o,open_n7680}),
    .b({_al_u1965_o,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .d({open_n7684,_al_u1965_o}),
    .sr(rst_pad),
    .q({open_n7702,\t/a/ID_rs2$1$_placeOpt_2 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_20  (
    .a({open_n7703,\t/a/if_id/n9 }),
    .b({_al_u1965_o,_al_u1965_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,open_n7707}),
    .sr(rst_pad),
    .q({open_n7725,\t/a/ID_rs2$1$_placeOpt_20 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_21  (
    .a({open_n7726,_al_u1965_o}),
    .c({_al_u1950_o,open_n7729}),
    .clk(clock_pad),
    .d({_al_u1965_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7748,\t/a/ID_rs2$1$_placeOpt_21 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0011000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_3  (
    .a({open_n7749,_al_u1965_o}),
    .b({_al_u1965_o,\t/a/if_id/n9 }),
    .c({_al_u1950_o,open_n7750}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n7771,\t/a/ID_rs2$1$_placeOpt_3 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0100010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_4  (
    .a({_al_u1965_o,_al_u1965_o}),
    .b({_al_u1950_o,open_n7772}),
    .clk(clock_pad),
    .d({open_n7776,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7794,\t/a/ID_rs2$1$_placeOpt_4 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B)"),
    //.LUT1("(~C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000011),
    .INIT_LUT1(16'b0000110000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_5  (
    .b({_al_u1950_o,\t/a/if_id/n9 }),
    .c({_al_u1965_o,_al_u1965_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n7817,\t/a/ID_rs2$1$_placeOpt_5 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~A*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0100010001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_6  (
    .a({_al_u1965_o,_al_u1965_o}),
    .b({_al_u1950_o,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n7840,\t/a/ID_rs2$1$_placeOpt_6 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_7  (
    .a({open_n7841,\t/a/if_id/n9 }),
    .b({_al_u1965_o,_al_u1965_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,open_n7845}),
    .sr(rst_pad),
    .q({open_n7863,\t/a/ID_rs2$1$_placeOpt_7 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_8  (
    .a({_al_u1965_o,\t/a/if_id/n9 }),
    .c({_al_u1950_o,_al_u1965_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n7886,\t/a/ID_rs2$1$_placeOpt_8 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1_placeOpt_9  (
    .a({_al_u1965_o,_al_u1965_o}),
    .c({_al_u1950_o,open_n7889}),
    .clk(clock_pad),
    .d({open_n7891,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n7909,\t/a/ID_rs2$1$_placeOpt_9 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(D*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1967|t/a/id_ex/reg3_b3  (
    .a({open_n7910,\t/a/aluin/sel1_b23/B9 }),
    .b({\t/a/MEM_rd [3],_al_u2007_o}),
    .c({open_n7911,_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_rs2 [3],\t/a/EX_rs2 [3]}),
    .mi({open_n7923,\t/a/ID_rs2$3$_placeOpt_3 }),
    .sr(rst_pad),
    .f({_al_u1967_o,\t/a/EX_B [23]}),
    .q({open_n7927,\t/a/EX_rs2 [3]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*A)"),
    //.LUT1("(B*D)"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b1100110000000000),
    .MODE("LOGIC"))
    \_al_u1972|_al_u1978  (
    .a({open_n7928,\t/a/n29 }),
    .b({\t/a/n24_lutinv ,open_n7929}),
    .d({_al_u1798_o,\t/a/n24_lutinv }),
    .f({\t/a/alu_B_select [0],\t/a/alu_B_select [1]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1973|t/a/id_ex/reg3_b0  (
    .a({open_n7952,\t/a/aluin/n12_lutinv }),
    .b({\t/a/WB_rd [0],_al_u1984_o}),
    .c({open_n7953,\t/a/EX_rs2 [0]}),
    .clk(clock_pad),
    .d({\t/a/EX_rs2 [0],\t/a/EX_rd [0]}),
    .mi({open_n7965,\t/a/ID_rs2$0$_placeOpt_21 }),
    .sr(rst_pad),
    .f({_al_u1973_o,_al_u2076_o}),
    .q({open_n7969,\t/a/EX_rs2 [0]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0@C)*~(D*~B))"),
    //.LUT1("(~A*~(1@C)*~(B*~D))"),
    .INIT_LUT0(16'b0000010000000101),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1974 (
    .a({_al_u1973_o,_al_u1973_o}),
    .b({\t/a/WB_rd [1],\t/a/EX_rs2 [1]}),
    .c({\t/a/EX_rs2 [3],\t/a/EX_rs2 [3]}),
    .d({\t/a/EX_rs2 [1],\t/a/WB_rd [1]}),
    .mi({open_n7982,\t/a/WB_rd [3]}),
    .fx({open_n7987,_al_u1974_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(~D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1975|t/a/id_ex/reg3_b1  (
    .a({open_n7990,\t/a/aluin/sel1_b21/B9 }),
    .b({open_n7991,_al_u2007_o}),
    .c({\t/a/EX_rs2 [1],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/WB_rd [1],\t/a/EX_rs2 [1]}),
    .mi({open_n8003,\t/a/ID_rs2$1$_placeOpt_15 }),
    .sr(rst_pad),
    .f({_al_u1975_o,\t/a/EX_B [21]}),
    .q({open_n8007,\t/a/EX_rs2 [1]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(A*B*C*~(0@D))"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(A*B*C*~(1@D))"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1977|_al_u1976  (
    .a({_al_u1976_o,_al_u1975_o}),
    .b({_al_u1974_o,\t/a/EX_rs2 [0]}),
    .c({\t/a/n19 ,\t/a/EX_rs2 [4]}),
    .d({\t/a/EX_rs2 [2],\t/a/WB_rd [0]}),
    .e({\t/a/WB_rd [2],\t/a/WB_rd [4]}),
    .f({\t/a/n29 ,_al_u1976_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~D*~C*~B+A*~D*~C*~B+A*~D*C*~B+~A*~D*~C*B+A*~D*~C*B+A*~D*C*B"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C"),
    //.LUTG0("~A*~D*~C*~B+~A*~D*~C*B"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000010101111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000000000000101),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1983|_al_u491  (
    .a({open_n8030,\t/a/ID_rs1$0$_placeOpt_20 }),
    .c({open_n8033,\t/a/regfile/regfile$4$ [31]}),
    .d({\t/a/aluin/n12_lutinv ,\t/a/ID_rs1$1$_placeOpt_20 }),
    .e({\t/a/aluin/n11_lutinv ,\t/a/regfile/regfile$5$ [31]}),
    .f({_al_u1983_o,_al_u491_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("B*~C*A*D+B*C*A*D"),
    //.LUTF1("0"),
    //.LUTG0("~B*~C*A*~D+B*~C*A*~D+~B*C*A*~D+B*C*A*~D+~B*~C*A*D+B*~C*A*D+~B*C*A*D+B*C*A*D"),
    //.LUTG1("~C*~A*~B*~D+C*~A*~B*~D+~C*A*~B*~D+C*A*~B*~D+~C*~A*~B*D+C*~A*~B*D+~C*A*~B*D+C*A*~B*D+~C*~A*B*D+~C*A*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101010),
    .INIT_LUTG1(16'b0011111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1985|t/a/ex_mem/reg3_b0  (
    .a({open_n8056,\t/a/EX_fun3 [0]}),
    .b({_al_u1984_o,_al_u1984_o}),
    .c({\t/a/EX_fun3 [1],open_n8057}),
    .clk(clock_pad),
    .d({\t/a/EX_fun3 [0],\t/a/EX_op [4]}),
    .e({_al_u1983_o,\t/a/aluin/n10_lutinv }),
    .mi({open_n8060,\t/a/EX_fun3 [0]}),
    .sr(rst_pad),
    .f({_al_u1985_o,\t/a/EX_operation [0]}),
    .q({open_n8075,\t/a/MEM_fun3 [0]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*B*A*~D+C*B*A*~D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("0"),
    //.LUTG0("~C*B*A*~D+C*B*A*~D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*C*D+B*~A*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010001000),
    .INIT_LUTG1(16'b0101000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1985|t/a/ex_mem/reg3_b0_placeOpt_1  (
    .a(\t/a/EX_fun3 [1:0]),
    .b({open_n8076,\t/a/aluin/n10_lutinv }),
    .c({\t/a/EX_fun3 [0],open_n8077}),
    .clk(clock_pad),
    .d({_al_u1984_o,\t/a/EX_op [4]}),
    .e({_al_u1983_o,_al_u1984_o}),
    .mi({open_n8080,\t/a/EX_fun3 [0]}),
    .sr(rst_pad),
    .f({open_n8092,\t/a/EX_operation$0$_lutinv_placeOpt_1 }));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*A*~C+D*B*A*~C+~D*B*A*C+D*B*A*C"),
    //.LUTF1("0"),
    //.LUTG0("D*~B*A*~C+~D*B*A*~C+D*B*A*~C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTG1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*C*D+B*~A*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010001000),
    .INIT_LUTG1(16'b0101000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1985|t/a/ex_mem/reg3_b0_placeOpt_2  (
    .a(\t/a/EX_fun3 [1:0]),
    .b({open_n8098,\t/a/aluin/n10_lutinv }),
    .c({\t/a/EX_fun3 [0],open_n8099}),
    .clk(clock_pad),
    .d({_al_u1984_o,_al_u1984_o}),
    .e({_al_u1983_o,\t/a/EX_op [4]}),
    .mi({open_n8102,\t/a/EX_fun3 [0]}),
    .sr(rst_pad),
    .f({open_n8114,\t/a/EX_operation$0$_lutinv_placeOpt_2 }));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*C*~A+D*B*C*~A+~D*B*C*A+D*B*C*A"),
    //.LUTF1("0"),
    //.LUTG0("D*~B*C*~A+~D*B*C*~A+D*B*C*~A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*~C*D+B*~A*~C*D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+~B*A*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000011000000),
    .INIT_LUTG1(16'b0011111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1985|t/a/ex_mem/reg3_b0_placeOpt_3  (
    .b({\t/a/EX_fun3 [1],\t/a/aluin/n10_lutinv }),
    .c({_al_u1984_o,\t/a/EX_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/EX_fun3 [0],_al_u1984_o}),
    .e({_al_u1983_o,\t/a/EX_op [4]}),
    .mi({open_n8124,\t/a/EX_fun3 [0]}),
    .sr(rst_pad),
    .f({open_n8136,\t/a/EX_operation$0$_lutinv_placeOpt_3 }));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~B*~(D*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(~B*~(D*A)))"),
    //.LUTG1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*C*D+B*~A*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110000011000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1110000011000000),
    .INIT_LUTG1(16'b0101000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1985|t/a/ex_mem/reg3_b0_placeOpt_4  (
    .a({\t/a/EX_fun3 [1],_al_u1984_o}),
    .b({open_n8142,\t/a/aluin/n10_lutinv }),
    .c({\t/a/EX_fun3 [0],\t/a/EX_fun3 [0]}),
    .clk(clock_pad),
    .d({_al_u1984_o,\t/a/EX_op [4]}),
    .e({_al_u1983_o,open_n8144}),
    .mi({open_n8146,\t/a/EX_fun3 [0]}),
    .sr(rst_pad),
    .f({open_n8158,\t/a/EX_operation$0$_lutinv_placeOpt_4 }));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("A*~C*~B*~D+A*C*~B*~D+A*~C*B*~D+A*C*B*~D+A*~C*B*D+A*C*B*D"),
    //.LUTG0("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("A*~C*~B*~D+A*C*~B*~D+A*~C*B*~D+A*C*B*~D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1000100010101010),
    .INIT_LUTG0(16'b1110111011001100),
    .INIT_LUTG1(16'b0000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1985|t/a/ex_mem/reg3_b0_placeOpt_5  (
    .a({_al_u1983_o,_al_u1984_o}),
    .b({\t/a/EX_fun3 [0],\t/a/aluin/n10_lutinv }),
    .clk(clock_pad),
    .d({_al_u1984_o,\t/a/EX_op [4]}),
    .e(\t/a/EX_fun3 [1:0]),
    .mi({open_n8168,\t/a/EX_fun3 [0]}),
    .sr(rst_pad),
    .f({open_n8180,\t/a/EX_operation$0$_lutinv_placeOpt_5 }));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~D*(B@A)))"),
    //.LUT1("~(~B*~(D*~A))"),
    .INIT_LUT0(16'b1111000010010000),
    .INIT_LUT1(16'b1101110111001100),
    .MODE("LOGIC"))
    \_al_u1986|_al_u2495  (
    .a({_al_u1985_o,\t/a/EX_A [9]}),
    .b({\t/a/aluin/sel1_b9/B9 ,\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o }),
    .c({open_n8186,_al_u2431_o}),
    .d({\t/a/EX_fun7 [4],\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .f({\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ,_al_u2495_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b0101000000000000),
    .INIT_LUTG1(16'b1111111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1989|t/a/regfile/reg0_b168  (
    .a({open_n8207,_al_u1987_o}),
    .b({_al_u1985_o,open_n8208}),
    .c({open_n8209,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b8/B9 ,\t/a/reg_writedat [8]}),
    .e({\t/a/EX_fun7 [3],\t/a/alu_B_select [1]}),
    .mi({open_n8211,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b8/B9 }),
    .q({open_n8226,\t/a/regfile/regfile$5$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("~C*~A*~B*~D+~C*~A*B*~D+~C*~A*~B*D+~C*A*~B*D+~C*~A*B*D+~C*A*B*D"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b0000111100000101),
    .INIT_LUTG1(16'b1111111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1992|t/a/regfile/reg0_b167  (
    .a({open_n8227,\t/a/alu_B_select [1]}),
    .c({_al_u1985_o,_al_u1990_o}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b7/B9 ,\t/a/reg_writedat [7]}),
    .e({\t/a/EX_fun7 [2],\t/a/aluin/n10_lutinv }),
    .mi({open_n8231,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/B9 }),
    .q({open_n8246,\t/a/regfile/regfile$5$ [7]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~A*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1011101110101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1995|t/a/regfile/reg0_b166  (
    .a({\t/a/aluin/sel1_b6/B9 ,_al_u1993_o}),
    .b({_al_u1985_o,\t/a/alu_B_select [1]}),
    .c({open_n8247,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [1],\t/a/reg_writedat [6]}),
    .mi({open_n8258,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b6/B9 }),
    .q({open_n8262,\t/a/regfile/regfile$5$ [6]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~A*~(B*~C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1010111010101110),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1998|t/a/regfile/reg0_b165  (
    .a({\t/a/aluin/sel1_b5/B9 ,_al_u1996_o}),
    .b({\t/a/EX_fun7 [0],\t/a/alu_B_select [1]}),
    .c({_al_u1985_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({open_n8263,\t/a/reg_writedat [5]}),
    .mi({open_n8274,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b5/B9 }),
    .q({open_n8278,\t/a/regfile/regfile$5$ [5]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~D*B*~A+~C*D*B*~A+~C*~D*B*A+~C*D*B*A"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~C*~D*B*A+~C*D*B*A"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110000001100),
    .INIT_LUTF1(16'b1111111110101010),
    .INIT_LUTG0(16'b0000100000001000),
    .INIT_LUTG1(16'b1111101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2004|t/a/regfile/reg0_b159  (
    .a({\t/a/aluin/sel1_b31/B9 ,\t/a/reg_writedat [31]}),
    .b({open_n8279,\t/a/aluin/n10_lutinv }),
    .c({_al_u1803_o,_al_u2002_o}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [6],open_n8280}),
    .e({_al_u1983_o,\t/a/alu_B_select [1]}),
    .mi({open_n8282,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [31],\t/a/aluin/sel1_b31/B9 }),
    .q({open_n8297,\t/a/regfile/regfile$4$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*C)"),
    //.LUTF1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(B*C)"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011000000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b1100000011000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2007|t/a/id_ex/reg2_b6  (
    .b({open_n8300,\t/a/ID_fun7 [6]}),
    .c({open_n8301,\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [6],open_n8303}),
    .e({_al_u1983_o,open_n8304}),
    .mi({open_n8306,\t/a/ID_fun7 [6]}),
    .sr(rst_pad),
    .f({_al_u2007_o,\t/a/condition/sel0_b12/B1 }),
    .q({open_n8321,\t/a/EX_fun7 [6]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111111111001100),
    .INIT_LUTG0(16'b0101010100010001),
    .INIT_LUTG1(16'b1111111111101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2008|t/a/regfile/reg0_b158  (
    .a({\t/a/EX_fun7 [5],_al_u2005_o}),
    .b({_al_u2007_o,\t/a/alu_B_select [1]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b30/B9 ,\t/a/reg_writedat [30]}),
    .e({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .mi({open_n8325,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [30],\t/a/aluin/sel1_b30/B9 }),
    .q({open_n8340,\t/a/regfile/regfile$4$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111011101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2014|t/a/regfile/reg0_b157  (
    .a({\t/a/aluin/sel1_b29/B9 ,_al_u2012_o}),
    .b({_al_u2007_o,\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [4],\t/a/reg_writedat [29]}),
    .mi({open_n8351,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [29],\t/a/aluin/sel1_b29/B9 }),
    .q({open_n8355,\t/a/regfile/regfile$4$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111011101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2017|t/a/regfile/reg0_b156  (
    .a({\t/a/aluin/sel1_b28/B9 ,_al_u2015_o}),
    .b({_al_u2007_o,\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [3],\t/a/reg_writedat [28]}),
    .mi({open_n8366,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [28],\t/a/aluin/sel1_b28/B9 }),
    .q({open_n8370,\t/a/regfile/regfile$4$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("A*~C*~B*~D+A*C*~B*~D+A*~C*B*~D+A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("A*~C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010000),
    .INIT_LUTF1(16'b1111111110101010),
    .INIT_LUTG0(16'b0101000000000000),
    .INIT_LUTG1(16'b1111111111101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2020|t/a/regfile/reg0_b155  (
    .a({\t/a/aluin/sel1_b27/B9 ,_al_u2018_o}),
    .b({_al_u1803_o,open_n8371}),
    .c({open_n8372,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2007_o,\t/a/reg_writedat [27]}),
    .e({\t/a/EX_fun7 [2],\t/a/alu_B_select [1]}),
    .mi({open_n8374,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [27],\t/a/aluin/sel1_b27/B9 }),
    .q({open_n8389,\t/a/regfile/regfile$4$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("A*~D*~B*~C+~A*D*~B*~C+A*D*~B*~C+A*~D*B*~C+~A*D*B*~C+A*D*B*~C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTG0("~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("A*~D*~B*~C+~A*D*~B*~C+A*D*~B*~C+~A*~D*B*~C+A*~D*B*~C+~A*D*B*~C+A*D*B*~C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010000),
    .INIT_LUTF1(16'b1111111110101010),
    .INIT_LUTG0(16'b0101000000000000),
    .INIT_LUTG1(16'b1111111111101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2023|t/a/regfile/reg0_b154  (
    .a({\t/a/aluin/sel1_b26/B9 ,_al_u2021_o}),
    .b({_al_u1803_o,open_n8390}),
    .c({open_n8391,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2007_o,\t/a/reg_writedat [26]}),
    .e({\t/a/EX_fun7 [1],\t/a/alu_B_select [1]}),
    .mi({open_n8393,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [26],\t/a/aluin/sel1_b26/B9 }),
    .q({open_n8408,\t/a/regfile/regfile$4$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~D*~A*~(B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111111101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2026|t/a/regfile/reg0_b153  (
    .a({\t/a/aluin/sel1_b25/B9 ,_al_u2024_o}),
    .b({\t/a/EX_fun7 [0],\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2007_o,\t/a/reg_writedat [25]}),
    .mi({open_n8419,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [25],\t/a/aluin/sel1_b25/B9 }),
    .q({open_n8423,\t/a/regfile/regfile$4$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111011101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2041|t/a/regfile/reg0_b148  (
    .a({\t/a/aluin/sel1_b20/B9 ,_al_u2039_o}),
    .b({_al_u2007_o,\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_rs2 [0],\t/a/reg_writedat [20]}),
    .mi({open_n8434,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [20],\t/a/aluin/sel1_b20/B9 }),
    .q({open_n8438,\t/a/regfile/regfile$4$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~D*(B@A)))"),
    //.LUT1("~(~B*~D*~(A*C))"),
    .INIT_LUT0(16'b1111000010010000),
    .INIT_LUT1(16'b1111111111101100),
    .MODE("LOGIC"))
    \_al_u2059|_al_u2445  (
    .a({\t/a/EX_fun3 [2],\t/a/EX_A [14]}),
    .b({_al_u2007_o,\t/a/EX_B [14]}),
    .c({_al_u1803_o,_al_u2431_o}),
    .d({\t/a/aluin/sel1_b14/B9 ,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .f({\t/a/EX_B [14],_al_u2445_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*B)"),
    //.LUT1("~(~B*~A*~(C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000100010001000),
    .INIT_LUT1(16'b1111111011101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2062|t/a/ex_mem/reg3_b1  (
    .a({\t/a/aluin/sel1_b13/B9 ,\t/a/EX_fun3 [1]}),
    .b({_al_u2007_o,\t/a/EX_operation [2]}),
    .c({\t/a/EX_fun3 [1],open_n8459}),
    .clk(clock_pad),
    .d({_al_u1803_o,open_n8461}),
    .mi({open_n8472,\t/a/EX_fun3 [1]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [13],_al_u2169_o}),
    .q({open_n8476,\t/a/MEM_fun3 [1]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*B*~D+~A*C*B*~D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTF1("A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("A*~C*B*~D+A*C*B*~D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG1("A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .INIT_LUTF0(16'b1100110001000100),
    .INIT_LUTF1(16'b1111101011111010),
    .INIT_LUTG0(16'b1100110010001000),
    .INIT_LUTG1(16'b1111111111111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2065|_al_u2465  (
    .a({\t/a/aluin/sel1_b12/B9 ,\t/a/EX_A [12]}),
    .b({open_n8477,_al_u2431_o}),
    .c({_al_u2007_o,open_n8478}),
    .d({_al_u1803_o,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .e({\t/a/EX_fun3 [0],\t/a/EX_B [12]}),
    .f({\t/a/EX_B [12],_al_u2465_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~A*B*~D+C*~A*B*~D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("~C*A*B*~D+C*A*B*~D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1100110001000100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1100110010001000),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2068|_al_u2475  (
    .a({open_n8501,\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o }),
    .b({open_n8502,_al_u2431_o}),
    .c({\t/a/EX_fun7 [6],open_n8503}),
    .d({_al_u1985_o,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .e({\t/a/aluin/sel1_b11/B9 ,\t/a/EX_A [11]}),
    .f({\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o ,_al_u2475_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~A*D*~C*~B+A*D*~C*~B+~A*D*C*~B+A*D*C*~B+~A*D*~C*B+A*D*~C*B+~A*D*C*B+A*D*C*B"),
    //.LUTG0("~C*~B*~A*~D+~C*~B*A*~D+~C*~B*~A*D+~C*B*~A*D+~C*~B*A*D+~C*B*A*D"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+~A*D*~C*B+A*D*~C*B+~A*D*C*B+A*D*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b0000111100000011),
    .INIT_LUTG1(16'b1111111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2071|t/a/regfile/reg0_b106  (
    .b({_al_u1985_o,\t/a/alu_B_select [1]}),
    .c({open_n8528,_al_u2069_o}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b10/B9 ,\t/a/reg_writedat [10]}),
    .e({\t/a/EX_fun7 [5],\t/a/aluin/n10_lutinv }),
    .mi({open_n8530,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b10/B9 }),
    .q({open_n8545,\t/a/regfile/regfile$3$ [10]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~A*~(~0*B)))"),
    //.LUT1("~(C*~(D*~A*~(~1*B)))"),
    .INIT_LUT0(16'b0001111100001111),
    .INIT_LUT1(16'b0101111100001111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2077 (
    .a({_al_u2075_o,_al_u2075_o}),
    .b({\t/a/alu_B_select [1],\t/a/alu_B_select [1]}),
    .c({_al_u2076_o,_al_u2076_o}),
    .d({\t/a/aluin/n10_lutinv ,\t/a/aluin/n10_lutinv }),
    .mi({open_n8558,\t/a/reg_writedat [0]}),
    .fx({open_n8563,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1011100000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2078|t/a/if_id/reg1_b6  (
    .a({i_data[31],\t/a/if_id/n9 }),
    .b({\t/busarbitration/n3_placeOpt_3 ,\t/busarbitration/n3_placeOpt_3 }),
    .c({\t/busarbitration/instruction [31],\t/busarbitration/instruction [31]}),
    .clk(clock_pad),
    .d({_al_u1950_o,i_data[31]}),
    .sr(rst_pad),
    .f({_al_u2078_o,open_n8579}),
    .q({open_n8583,\t/a/ID_fun7 [6]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~((0*D))*~(A)+(C*B)*(0*D)*~(A)+~((C*B))*(0*D)*A+(C*B)*(0*D)*A)"),
    //.LUTF1("~((~C*~A)*~((~0*~B))*~(D)+(~C*~A)*(~0*~B)*~(D)+~((~C*~A))*(~0*~B)*D+(~C*~A)*(~0*~B)*D)"),
    //.LUTG0("~((C*B)*~((1*D))*~(A)+(C*B)*(1*D)*~(A)+~((C*B))*(1*D)*A+(C*B)*(1*D)*A)"),
    //.LUTG1("~((~C*~A)*~((~1*~B))*~(D)+(~C*~A)*(~1*~B)*~(D)+~((~C*~A))*(~1*~B)*D+(~C*~A)*(~1*~B)*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011111110111111),
    .INIT_LUTF1(16'b1100110011111010),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b1111111111111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2079|_al_u1944  (
    .a({\t/busarbitration/instruction [5],\t/busarbitration/n3_placeOpt_2 }),
    .b({i_data[6],\t/busarbitration/instruction [5]}),
    .c({\t/busarbitration/instruction [6],\t/busarbitration/instruction [6]}),
    .clk(clock_pad),
    .d({\t/busarbitration/n3_placeOpt_2 ,i_data[6]}),
    .e({i_data[5],i_data[5]}),
    .mi({i_data[6],i_data[6]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({\t/a/unconditional/eq1/or_xor_i0$5$_i1$5$_o_o_lutinv ,_al_u1944_o}),
    .q({\trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*C*~B*~A)"),
    //.LUT1("(~1*~D*C*~B*~A)"),
    .INIT_LUT0(16'b0000000000010000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2080 (
    .a({_al_u1948_o,_al_u1948_o}),
    .b({\t/instruction$2$_neg_lutinv ,\t/instruction$2$_neg_lutinv }),
    .c({\t/instruction$3$_neg_lutinv ,\t/instruction$3$_neg_lutinv }),
    .d({\t/instruction$4$_neg_lutinv ,\t/instruction$4$_neg_lutinv }),
    .mi({open_n8612,\t/a/unconditional/eq1/or_xor_i0$5$_i1$5$_o_o_lutinv }),
    .fx({open_n8617,_al_u2080_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUT1("~(~A*~(B*(C*~(1)*~(D)+C*1*~(D)+~(C)*1*D+C*1*D)))"),
    .INIT_LUT0(16'b1010111010101010),
    .INIT_LUT1(16'b1110111011101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2081 (
    .a({_al_u2078_o,_al_u2078_o}),
    .b({_al_u2080_o,_al_u2080_o}),
    .c({\t/busarbitration/instruction [30],\t/busarbitration/n3_placeOpt_3 }),
    .d({\t/busarbitration/n3_placeOpt_3 ,\t/busarbitration/instruction [30]}),
    .mi({open_n8632,i_data[30]}),
    .fx({open_n8637,\t/a/IF_skip_addr [30]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUT1("~(~A*~(B*(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111010101010),
    .INIT_LUT1(16'b1110111011101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    _al_u2082 (
    .a({_al_u2078_o,_al_u2078_o}),
    .b({_al_u2080_o,_al_u2080_o}),
    .c({\t/busarbitration/n3_placeOpt_4 ,\t/busarbitration/n3_placeOpt_4 }),
    .clk(clock_pad),
    .d({\t/busarbitration/instruction [29],\t/busarbitration/instruction [29]}),
    .mi({i_data[29],i_data[29]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .fx({open_n8654,\t/a/IF_skip_addr [29]}),
    .q({\trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/ctl_this ,open_n8655}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUT1("~(~A*~(B*(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .INIT_LUT0(16'b1010111010101010),
    .INIT_LUT1(16'b1110111011101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2085 (
    .a({_al_u2078_o,_al_u2078_o}),
    .b({_al_u2080_o,_al_u2080_o}),
    .c({\t/busarbitration/n3_placeOpt_3 ,\t/busarbitration/n3_placeOpt_3 }),
    .d({\t/busarbitration/instruction [26],\t/busarbitration/instruction [26]}),
    .mi({open_n8668,i_data[26]}),
    .fx({open_n8673,\t/a/IF_skip_addr [26]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUT1("~(~A*~(B*(C*~(1)*~(D)+C*1*~(D)+~(C)*1*D+C*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111010101010),
    .INIT_LUT1(16'b1110111011101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    _al_u2086 (
    .a({_al_u2078_o,_al_u2078_o}),
    .b({_al_u2080_o,_al_u2080_o}),
    .c({\t/busarbitration/instruction [25],\t/busarbitration/n3_placeOpt_3 }),
    .clk(clock_pad),
    .d({\t/busarbitration/n3_placeOpt_3 ,\t/busarbitration/instruction [25]}),
    .mi({i_data[25],i_data[25]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .fx({open_n8690,\t/a/IF_skip_addr [25]}),
    .q({\trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/level_0_r ,open_n8691}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(~C*B))"),
    //.LUTF1("D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("~(~D*~(~C*B))"),
    //.LUTG1("D*~B*~C*~A+D*B*~C*~A+D*~B*C*~A+D*B*C*~A+D*~B*~C*A+D*B*~C*A+D*~B*C*A+D*B*C*A"),
    .INIT_LUTF0(16'b1111111100001100),
    .INIT_LUTF1(16'b1111111111001100),
    .INIT_LUTG0(16'b1111111100001100),
    .INIT_LUTG1(16'b1111111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2087|_al_u2089  (
    .b({_al_u2080_o,_al_u2080_o}),
    .c({open_n8694,_al_u1960_o}),
    .d({_al_u2078_o,_al_u2078_o}),
    .e({_al_u1956_o,open_n8697}),
    .f({\t/a/IF_skip_addr [24],\t/a/IF_skip_addr [22]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    //.LUT1("~(~C*~(~A*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010100110011),
    .INIT_LUT1(16'b1111010011110100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2088|_al_u1958  (
    .a({_al_u1958_o,i_data[23]}),
    .b({_al_u2080_o,\t/busarbitration/instruction [23]}),
    .c({_al_u2078_o,open_n8718}),
    .clk(clock_pad),
    .d({open_n8720,\t/busarbitration/n3_placeOpt_5 }),
    .mi({open_n8731,i_data[23]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({\t/a/IF_skip_addr [23],_al_u1958_o}),
    .q({open_n8735,\trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/ctl_this }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D)"),
    //.LUTF1("~A*B*~C*~D+~A*B*C*~D+~A*B*~C*D+~A*B*C*D"),
    //.LUTG0("~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111101010101),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b0000111101010101),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2090|_al_u1965  (
    .a({_al_u1965_o,\t/busarbitration/instruction [21]}),
    .b({_al_u2080_o,open_n8736}),
    .c({open_n8737,i_data[21]}),
    .clk(clock_pad),
    .d({open_n8739,\t/busarbitration/n3_placeOpt_2 }),
    .e({_al_u2078_o,open_n8740}),
    .mi({i_data[21],i_data[21]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({\t/a/IF_skip_addr [21],_al_u1965_o}),
    .q({\trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*A*~C*~D+B*A*~C*~D+~B*A*C*~D+B*A*C*~D"),
    //.LUTF1("~D*~B*~C*~A+~D*~B*~C*A"),
    //.LUTG0("~B*A*~C*~D+B*A*~C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG1("0"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1111111110101010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2095|t/a/if_id/reg5_b22  (
    .a({open_n8756,\t/a/MEM_aludat [22]}),
    .b({addr[21],open_n8757}),
    .c({addr[20],open_n8758}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[22],\t/busarbitration/n3_placeOpt_4 }),
    .e({addr[2],\t/memstraddress [22]}),
    .mi({open_n8760,\t/memstraddress [22]}),
    .sr(rst_pad),
    .f({_al_u2095_o,addr[22]}),
    .q({open_n8775,\t/a/ID_memstraddr [22]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*~C*~D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011001100),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2096|t/a/if_id/reg5_b19  (
    .a({addr[16],open_n8776}),
    .b({addr[19],\t/a/MEM_aludat [19]}),
    .c({addr[18],\t/memstraddress [19]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[17],open_n8777}),
    .e({_al_u2095_o,\t/busarbitration/n3_placeOpt_1 }),
    .mi({open_n8779,\t/memstraddress [19]}),
    .sr(rst_pad),
    .f({_al_u2096_o,addr[19]}),
    .q({open_n8794,\t/a/ID_memstraddr [19]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*A*B)"),
    //.LUTF1("(D*~C)"),
    //.LUTG0("(1*D*C*A*B)"),
    //.LUTG1("(D*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2097|_al_u2101  (
    .a({open_n8795,_al_u2097_o}),
    .b({open_n8796,_al_u2096_o}),
    .c({addr[11],_al_u2098_o}),
    .clk(clock_pad),
    .d({addr[10],_al_u2099_o}),
    .e({open_n8798,_al_u2100_o}),
    .mi({addr[11],addr[11]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u2097_o,_al_u2101_o}),
    .q({\trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*A)"),
    //.LUT1("(~D*C)"),
    .INIT_LUT0(16'b1010000010100000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u2098|_al_u1738  (
    .a({open_n8814,_al_u1735_o}),
    .c({addr[1],_al_u1737_o}),
    .d({addr[0],open_n8819}),
    .f({_al_u2098_o,\t/a/risk_jump/n35_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~B)"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B"),
    //.LUTG0("(~A*~B)"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001000100010001),
    .INIT_LUTF1(16'b0011001100110011),
    .INIT_LUTG0(16'b0001000100010001),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2099|_al_u2100  (
    .a({open_n8838,addr[12]}),
    .b(addr[14:13]),
    .clk(clock_pad),
    .e({addr[15],open_n8844}),
    .mi({addr[15],addr[15]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u2099_o,_al_u2100_o}),
    .q({\trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D"),
    //.LUTG0("(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    //.LUTG1("0"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011001100),
    .INIT_LUTF1(16'b0000000000000101),
    .INIT_LUTG0(16'b1010101011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2102|t/a/if_id/reg5_b31  (
    .a({addr[4],\t/memstraddress [31]}),
    .b({open_n8860,\t/a/MEM_aludat [31]}),
    .c({addr[31],open_n8861}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[30],\t/busarbitration/n3_placeOpt_4 }),
    .e({addr[5],open_n8862}),
    .mi({open_n8864,\t/memstraddress [31]}),
    .sr(rst_pad),
    .f({_al_u2102_o,addr[31]}),
    .q({open_n8879,\t/a/ID_memstraddr [31]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~D*~C+A*B*~D*~C+~A*B*D*~C+A*B*D*~C+~A*B*~D*C+A*B*~D*C+~A*B*D*C+A*B*D*C"),
    //.LUTF1("~A*B*~C*~D+~A*B*C*~D+~A*B*~C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG1("0"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011001100),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2103|t/a/if_id/reg5_b9  (
    .a({\t/a/MEM_aludat [9],open_n8880}),
    .b({memwrite_cs,\t/a/MEM_aludat [9]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({open_n8883,\t/memstraddress [9]}),
    .e({addr[8],\t/busarbitration/n3_placeOpt_5 }),
    .mi({open_n8885,\t/memstraddress [9]}),
    .sr(rst_pad),
    .f({_al_u2103_o,addr[9]}),
    .q({open_n8900,\t/a/ID_memstraddr [9]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    //.LUT1("(~D*~C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010110010101100),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2104|t/a/if_id/reg5_b7  (
    .a({_al_u2102_o,\t/memstraddress [7]}),
    .b({_al_u2103_o,\t/a/MEM_aludat [7]}),
    .c({addr[7],\t/busarbitration/n3_placeOpt_3 }),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[6],open_n8901}),
    .mi({open_n8912,\t/memstraddress [7]}),
    .sr(rst_pad),
    .f({_al_u2104_o,addr[7]}),
    .q({open_n8916,\t/a/ID_memstraddr [7]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~C*~A*~B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2105|t/a/if_id/reg5_b29  (
    .a({addr[29],open_n8917}),
    .b({addr[3],\t/a/MEM_aludat [29]}),
    .c({addr[28],\t/memstraddress [29]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[27],\t/busarbitration/n3_placeOpt_4 }),
    .mi({open_n8928,\t/memstraddress [29]}),
    .sr(rst_pad),
    .f({_al_u2105_o,addr[29]}),
    .q({open_n8932,\t/a/ID_memstraddr [29]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*C*~B*~D+A*C*~B*~D+~A*C*B*~D+A*C*B*~D+~A*C*~B*D+A*C*~B*D+~A*C*B*D+A*C*B*D"),
    //.LUTF1("(~B*~A)"),
    //.LUTG0("A*~C*~B*~D+A*C*~B*~D+A*~C*B*~D+A*C*B*~D+A*~C*~B*D+A*C*~B*D+A*~C*B*D+A*C*B*D"),
    //.LUTG1("(~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b1010101010101010),
    .INIT_LUTG1(16'b0001000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2106|t/a/if_id/reg5_b26  (
    .a({addr[26],\t/memstraddress [26]}),
    .b({addr[25],open_n8933}),
    .c({open_n8934,\t/a/MEM_aludat [26]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .e({open_n8937,\t/busarbitration/n3_placeOpt_4 }),
    .mi({open_n8939,\t/memstraddress [26]}),
    .sr(rst_pad),
    .f({_al_u2106_o,addr[26]}),
    .q({open_n8954,\t/a/ID_memstraddr [26]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUT1("(~C*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110010011100100),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2107|t/a/if_id/reg5_b24  (
    .a({addr[24],\t/busarbitration/n3_placeOpt_4 }),
    .b({open_n8955,\t/a/MEM_aludat [24]}),
    .c({addr[23],\t/memstraddress [24]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .mi({open_n8968,\t/memstraddress [24]}),
    .sr(rst_pad),
    .f({_al_u2107_o,addr[24]}),
    .q({open_n8972,\t/a/ID_memstraddr [24]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(0*D*C*B*A)"),
    //.LUT1("(1*D*C*B*A)"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2108 (
    .a({_al_u2101_o,_al_u2101_o}),
    .b({_al_u2104_o,_al_u2104_o}),
    .c({_al_u2105_o,_al_u2105_o}),
    .d({_al_u2106_o,_al_u2106_o}),
    .mi({open_n8985,_al_u2107_o}),
    .fx({open_n8990,n7}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*C*~D*B+A*C*D*B"),
    //.LUTF1("(~B*~C)"),
    //.LUTG0("A*~C*~D*~B+A*~C*D*~B+A*~C*~D*B+A*C*~D*B+A*~C*D*B+A*C*D*B"),
    //.LUTG1("(~B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000010000000),
    .INIT_LUTF1(16'b0000001100000011),
    .INIT_LUTG0(16'b1000101010001010),
    .INIT_LUTG1(16'b0000001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2109|_al_u1954  (
    .a({open_n8993,_al_u1950_o}),
    .b({_al_u2080_o,i_data[26]}),
    .c({_al_u1950_o,\t/busarbitration/n3_placeOpt_3 }),
    .clk(clock_pad),
    .e({open_n8997,\t/busarbitration/instruction [26]}),
    .mi({i_data[26],i_data[26]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u2109_o,\t/a/IF_skip_addr [6]}),
    .q({\trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111111111111),
    .INIT_LUTF1(16'b1111111100110011),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2111|_al_u2113  (
    .b({\t/busarbitration/instruction [19],open_n9015}),
    .c({open_n9016,i_data[18]}),
    .clk(clock_pad),
    .d({\t/busarbitration/n3_placeOpt_5 ,\t/busarbitration/n3_placeOpt_5 }),
    .e({i_data[19],\t/busarbitration/instruction [18]}),
    .mi({i_data[19],i_data[19]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({_al_u2111_o,_al_u2113_o}),
    .q({\trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~A)"),
    //.LUTF1("(~B*~D)"),
    //.LUTG0("(~B*~A)"),
    //.LUTG1("(~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001000100010001),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b0001000100010001),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2112|t/a/if_id/reg3_b4  (
    .a({open_n9033,\t/a/if_id/n9 }),
    .b({_al_u2111_o,_al_u2111_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,open_n9037}),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [19],open_n9054}),
    .q({open_n9058,\t/a/ID_rs1 [4]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2114|t/a/if_id/reg3_b3  (
    .b({_al_u2113_o,_al_u2113_o}),
    .c({_al_u2109_o,open_n9061}),
    .clk(clock_pad),
    .d({open_n9063,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [18],open_n9076}),
    .q({open_n9080,\t/a/ID_rs1 [3]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2114|t/a/if_id/reg3_b3_placeOpt_1  (
    .a({_al_u2113_o,_al_u2113_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9103,\t/a/ID_rs1$3$_placeOpt_1 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2114|t/a/if_id/reg3_b3_placeOpt_2  (
    .a({_al_u2109_o,open_n9104}),
    .c({_al_u2113_o,_al_u2113_o}),
    .clk(clock_pad),
    .d({open_n9108,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9126,\t/a/ID_rs1$3$_placeOpt_2 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B)"),
    //.LUT1("(~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000011),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2114|t/a/if_id/reg3_b3_placeOpt_3  (
    .a({_al_u2109_o,open_n9127}),
    .b({_al_u2113_o,\t/a/if_id/n9 }),
    .c({open_n9128,_al_u2113_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n9149,\t/a/ID_rs1$3$_placeOpt_3 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)"),
    //.LUT1("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001101010101),
    .INIT_LUT1(16'b0001101100011011),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2115|_al_u2119  (
    .a({\t/busarbitration/n3_placeOpt_5 ,\t/busarbitration/instruction [15]}),
    .b({\t/busarbitration/instruction [17],i_data[15]}),
    .c({i_data[17],open_n9150}),
    .clk(clock_pad),
    .d({open_n9152,\t/busarbitration/n3_placeOpt_5 }),
    .mi({i_data[17],i_data[17]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({_al_u2115_o,_al_u2119_o}),
    .q({\trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2  (
    .a({_al_u2109_o,open_n9166}),
    .c({_al_u2115_o,_al_u2115_o}),
    .clk(clock_pad),
    .d({open_n9170,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [17],open_n9183}),
    .q({open_n9187,\t/a/ID_rs1 [2]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2_placeOpt_1  (
    .b({_al_u2115_o,_al_u2115_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9210,\t/a/ID_rs1$2$_placeOpt_1 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~A*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2_placeOpt_10  (
    .a({_al_u2115_o,\t/a/if_id/n9 }),
    .b({open_n9211,_al_u2115_o}),
    .c({_al_u2109_o,open_n9212}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n9233,\t/a/ID_rs1$2$_placeOpt_10 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(~B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2_placeOpt_2  (
    .b({_al_u2115_o,\t/a/if_id/n9 }),
    .c({_al_u2109_o,open_n9236}),
    .clk(clock_pad),
    .d({open_n9238,_al_u2115_o}),
    .sr(rst_pad),
    .q({open_n9256,\t/a/ID_rs1$2$_placeOpt_2 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~A*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2_placeOpt_3  (
    .a({_al_u2115_o,open_n9257}),
    .b({_al_u2109_o,open_n9258}),
    .c({open_n9259,_al_u2115_o}),
    .clk(clock_pad),
    .d({open_n9261,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9279,\t/a/ID_rs1$2$_placeOpt_3 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A)"),
    //.LUT1("(~A*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2_placeOpt_4  (
    .a({_al_u2115_o,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .d({_al_u2109_o,_al_u2115_o}),
    .sr(rst_pad),
    .q({open_n9302,\t/a/ID_rs1$2$_placeOpt_4 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2_placeOpt_5  (
    .a({_al_u2109_o,open_n9303}),
    .c({_al_u2115_o,_al_u2115_o}),
    .clk(clock_pad),
    .d({open_n9307,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9325,\t/a/ID_rs1$2$_placeOpt_5 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~A*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2_placeOpt_6  (
    .a({_al_u2115_o,_al_u2115_o}),
    .b({open_n9326,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .d({_al_u2109_o,open_n9330}),
    .sr(rst_pad),
    .q({open_n9348,\t/a/ID_rs1$2$_placeOpt_6 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2_placeOpt_7  (
    .a({_al_u2109_o,open_n9349}),
    .c({_al_u2115_o,_al_u2115_o}),
    .clk(clock_pad),
    .d({open_n9353,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9371,\t/a/ID_rs1$2$_placeOpt_7 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2_placeOpt_8  (
    .b({_al_u2115_o,_al_u2115_o}),
    .c({_al_u2109_o,open_n9374}),
    .clk(clock_pad),
    .d({open_n9376,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9394,\t/a/ID_rs1$2$_placeOpt_8 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~A*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2_placeOpt_9  (
    .a({_al_u2115_o,_al_u2115_o}),
    .b({_al_u2109_o,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n9417,\t/a/ID_rs1$2$_placeOpt_9 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1  (
    .b({_al_u2117_o,_al_u2117_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [16],open_n9435}),
    .q({open_n9439,\t/a/ID_rs1 [1]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~A*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_1  (
    .a({_al_u2117_o,\t/a/if_id/n9 }),
    .b({open_n9440,_al_u2117_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,open_n9444}),
    .sr(rst_pad),
    .q({open_n9462,\t/a/ID_rs1$1$_placeOpt_1 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_10  (
    .a({_al_u2117_o,_al_u2117_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9485,\t/a/ID_rs1$1$_placeOpt_10 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~A*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_11  (
    .a({_al_u2117_o,_al_u2117_o}),
    .b({_al_u2109_o,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n9508,\t/a/ID_rs1$1$_placeOpt_11 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_12  (
    .c({_al_u2117_o,_al_u2117_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9531,\t/a/ID_rs1$1$_placeOpt_12 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_13  (
    .a({_al_u2117_o,_al_u2117_o}),
    .c({_al_u2109_o,open_n9534}),
    .clk(clock_pad),
    .d({open_n9536,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9554,\t/a/ID_rs1$1$_placeOpt_13 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_14  (
    .b({_al_u2109_o,open_n9557}),
    .c({_al_u2117_o,_al_u2117_o}),
    .clk(clock_pad),
    .d({open_n9559,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9577,\t/a/ID_rs1$1$_placeOpt_14 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(~B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_15  (
    .b({_al_u2117_o,\t/a/if_id/n9 }),
    .c({_al_u2109_o,open_n9580}),
    .clk(clock_pad),
    .d({open_n9582,_al_u2117_o}),
    .sr(rst_pad),
    .q({open_n9600,\t/a/ID_rs1$1$_placeOpt_15 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_16  (
    .c({_al_u2117_o,_al_u2117_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9623,\t/a/ID_rs1$1$_placeOpt_16 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B)"),
    //.LUT1("(~C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000011),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_17  (
    .a({_al_u2109_o,open_n9624}),
    .b({open_n9625,\t/a/if_id/n9 }),
    .c({_al_u2117_o,_al_u2117_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n9646,\t/a/ID_rs1$1$_placeOpt_17 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A)"),
    //.LUT1("(~C*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_18  (
    .a({open_n9647,\t/a/if_id/n9 }),
    .b({_al_u2109_o,open_n9648}),
    .c({_al_u2117_o,_al_u2117_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n9669,\t/a/ID_rs1$1$_placeOpt_18 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_19  (
    .a({_al_u2117_o,_al_u2117_o}),
    .b({_al_u2109_o,open_n9670}),
    .clk(clock_pad),
    .d({open_n9674,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9692,\t/a/ID_rs1$1$_placeOpt_19 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_2  (
    .a({open_n9693,\t/a/if_id/n9 }),
    .b({_al_u2117_o,_al_u2117_o}),
    .c({_al_u2109_o,open_n9694}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n9715,\t/a/ID_rs1$1$_placeOpt_2 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_20  (
    .b({_al_u2109_o,open_n9718}),
    .c({_al_u2117_o,_al_u2117_o}),
    .clk(clock_pad),
    .d({open_n9720,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9738,\t/a/ID_rs1$1$_placeOpt_20 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~A*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_21  (
    .a({_al_u2117_o,_al_u2117_o}),
    .b({open_n9739,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .d({_al_u2109_o,open_n9743}),
    .sr(rst_pad),
    .q({open_n9761,\t/a/ID_rs1$1$_placeOpt_21 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~A*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_3  (
    .a({_al_u2117_o,\t/a/if_id/n9 }),
    .b({open_n9762,_al_u2117_o}),
    .c({_al_u2109_o,open_n9763}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n9784,\t/a/ID_rs1$1$_placeOpt_3 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_4  (
    .a({open_n9785,\t/a/if_id/n9 }),
    .b({_al_u2117_o,_al_u2117_o}),
    .c({_al_u2109_o,open_n9786}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n9807,\t/a/ID_rs1$1$_placeOpt_4 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_5  (
    .a({_al_u2117_o,_al_u2117_o}),
    .b({_al_u2109_o,open_n9808}),
    .clk(clock_pad),
    .d({open_n9812,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9830,\t/a/ID_rs1$1$_placeOpt_5 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_6  (
    .a({_al_u2109_o,open_n9831}),
    .b({_al_u2117_o,_al_u2117_o}),
    .clk(clock_pad),
    .d({open_n9835,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9853,\t/a/ID_rs1$1$_placeOpt_6 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_7  (
    .a({open_n9854,_al_u2117_o}),
    .b({_al_u2117_o,\t/a/if_id/n9 }),
    .c({_al_u2109_o,open_n9855}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n9876,\t/a/ID_rs1$1$_placeOpt_7 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_8  (
    .a({_al_u2109_o,\t/a/if_id/n9 }),
    .b({_al_u2117_o,_al_u2117_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n9899,\t/a/ID_rs1$1$_placeOpt_8 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1_placeOpt_9  (
    .a({_al_u2117_o,_al_u2117_o}),
    .b({_al_u2109_o,open_n9900}),
    .clk(clock_pad),
    .d({open_n9904,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9922,\t/a/ID_rs1$1$_placeOpt_9 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0  (
    .b({_al_u2119_o,_al_u2119_o}),
    .c({_al_u2109_o,open_n9925}),
    .clk(clock_pad),
    .d({open_n9927,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [15],open_n9940}),
    .q({open_n9944,\t/a/ID_rs1 [0]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~D*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_1  (
    .b({open_n9947,_al_u2119_o}),
    .c({_al_u2109_o,open_n9948}),
    .clk(clock_pad),
    .d({_al_u2119_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9967,\t/a/ID_rs1$0$_placeOpt_1 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_10  (
    .b({_al_u2119_o,_al_u2119_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n9990,\t/a/ID_rs1$0$_placeOpt_10 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A)"),
    //.LUT1("(~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_11  (
    .a({_al_u2109_o,\t/a/if_id/n9 }),
    .b({_al_u2119_o,open_n9991}),
    .clk(clock_pad),
    .d({open_n9995,_al_u2119_o}),
    .sr(rst_pad),
    .q({open_n10013,\t/a/ID_rs1$0$_placeOpt_11 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A)"),
    //.LUT1("(~C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_12  (
    .a({_al_u2109_o,\t/a/if_id/n9 }),
    .c({_al_u2119_o,_al_u2119_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n10036,\t/a/ID_rs1$0$_placeOpt_12 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~B)"),
    //.LUT1("(~D*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_13  (
    .a({_al_u2109_o,open_n10037}),
    .b({open_n10038,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .d({_al_u2119_o,_al_u2119_o}),
    .sr(rst_pad),
    .q({open_n10059,\t/a/ID_rs1$0$_placeOpt_13 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000010100000101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_14  (
    .a({_al_u2109_o,open_n10060}),
    .c({_al_u2119_o,_al_u2119_o}),
    .clk(clock_pad),
    .d({open_n10064,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n10082,\t/a/ID_rs1$0$_placeOpt_14 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010100000101),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_15  (
    .a({open_n10083,\t/a/if_id/n9 }),
    .c({_al_u2119_o,_al_u2119_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,open_n10087}),
    .sr(rst_pad),
    .q({open_n10105,\t/a/ID_rs1$0$_placeOpt_15 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~D*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_16  (
    .a({_al_u2109_o,open_n10106}),
    .c({open_n10109,_al_u2119_o}),
    .clk(clock_pad),
    .d({_al_u2119_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n10128,\t/a/ID_rs1$0$_placeOpt_16 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A)"),
    //.LUT1("(~C*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_17  (
    .a({open_n10129,\t/a/if_id/n9 }),
    .b({_al_u2109_o,open_n10130}),
    .c({_al_u2119_o,open_n10131}),
    .clk(clock_pad),
    .d({open_n10133,_al_u2119_o}),
    .sr(rst_pad),
    .q({open_n10151,\t/a/ID_rs1$0$_placeOpt_17 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B)"),
    //.LUT1("(~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000011),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_18  (
    .a({_al_u2109_o,open_n10152}),
    .b({_al_u2119_o,\t/a/if_id/n9 }),
    .c({open_n10153,_al_u2119_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n10174,\t/a/ID_rs1$0$_placeOpt_18 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~B)"),
    //.LUT1("(~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001100000011),
    .INIT_LUT1(16'b0000000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_19  (
    .b({_al_u2119_o,\t/a/if_id/n9 }),
    .c({open_n10177,_al_u2119_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,open_n10179}),
    .sr(rst_pad),
    .q({open_n10197,\t/a/ID_rs1$0$_placeOpt_19 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A)"),
    //.LUT1("(~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_2  (
    .a({open_n10198,\t/a/if_id/n9 }),
    .b({_al_u2119_o,open_n10199}),
    .clk(clock_pad),
    .d({_al_u2109_o,_al_u2119_o}),
    .sr(rst_pad),
    .q({open_n10220,\t/a/ID_rs1$0$_placeOpt_2 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~A*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_20  (
    .a({_al_u2119_o,_al_u2119_o}),
    .b({open_n10221,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .d({_al_u2109_o,open_n10225}),
    .sr(rst_pad),
    .q({open_n10243,\t/a/ID_rs1$0$_placeOpt_20 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~A)"),
    //.LUT1("(~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_21  (
    .a({_al_u2109_o,\t/a/if_id/n9 }),
    .b({_al_u2119_o,_al_u2119_o}),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n10266,\t/a/ID_rs1$0$_placeOpt_21 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_3  (
    .b({_al_u2119_o,open_n10269}),
    .c({_al_u2109_o,_al_u2119_o}),
    .clk(clock_pad),
    .d({open_n10271,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n10289,\t/a/ID_rs1$0$_placeOpt_3 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A)"),
    //.LUT1("(~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_4  (
    .a({_al_u2109_o,\t/a/if_id/n9 }),
    .b({_al_u2119_o,open_n10290}),
    .clk(clock_pad),
    .d({open_n10294,_al_u2119_o}),
    .sr(rst_pad),
    .q({open_n10312,\t/a/ID_rs1$0$_placeOpt_4 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~D)"),
    //.LUT1("(~A*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000000001010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_5  (
    .a({_al_u2119_o,_al_u2119_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n10335,\t/a/ID_rs1$0$_placeOpt_5 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(~B*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b0000001100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_6  (
    .b({_al_u2119_o,_al_u2119_o}),
    .c({_al_u2109_o,open_n10338}),
    .clk(clock_pad),
    .d({open_n10340,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .q({open_n10358,\t/a/ID_rs1$0$_placeOpt_6 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A)"),
    //.LUT1("(~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_7  (
    .a({open_n10359,\t/a/if_id/n9 }),
    .b({_al_u2119_o,open_n10360}),
    .clk(clock_pad),
    .d({_al_u2109_o,_al_u2119_o}),
    .sr(rst_pad),
    .q({open_n10381,\t/a/ID_rs1$0$_placeOpt_7 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A)"),
    //.LUT1("(~D*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_8  (
    .a({open_n10382,\t/a/if_id/n9 }),
    .b({_al_u2109_o,open_n10383}),
    .clk(clock_pad),
    .d({_al_u2119_o,_al_u2119_o}),
    .sr(rst_pad),
    .q({open_n10404,\t/a/ID_rs1$0$_placeOpt_8 }));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~B)"),
    //.LUT1("(~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001000100010001),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0_placeOpt_9  (
    .a({_al_u2109_o,_al_u2119_o}),
    .b({_al_u2119_o,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .sr(rst_pad),
    .q({open_n10427,\t/a/ID_rs1$0$_placeOpt_9 }));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*A*~C+B*~D*A*~C+~B*D*~A*C+B*D*~A*C+~B*~D*A*C+B*~D*A*C+~B*D*A*C+B*D*A*C"),
    //.LUTF1("~A*D*~B*C+~A*D*B*C"),
    //.LUTG0("0"),
    //.LUTG1("~A*~D*~B*~C+~A*~D*B*~C+~A*~D*~B*C+~A*D*~B*C+~A*~D*B*C+~A*D*B*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000010101010),
    .INIT_LUTF1(16'b0101000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0101000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2121|t/a/if_id/reg0_b2  (
    .a({_al_u2109_o,\t/busarbitration/instruction [14]}),
    .c({i_data[14],i_data[14]}),
    .clk(clock_pad),
    .d({\t/busarbitration/n3_placeOpt_5 ,\t/busarbitration/n3_placeOpt_5 }),
    .e({\t/busarbitration/instruction [14],\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [14],open_n10445}),
    .q({open_n10449,\t/a/ID_fun3 [2]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0101010000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2122|t/a/if_id/reg0_b1  (
    .a({_al_u2109_o,\t/a/if_id/n9 }),
    .b({\t/busarbitration/n3_placeOpt_3 ,\t/busarbitration/n3_placeOpt_3 }),
    .c({\t/busarbitration/instruction [13],\t/busarbitration/instruction [13]}),
    .clk(clock_pad),
    .d({i_data[13],i_data[13]}),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [13],open_n10463}),
    .q({open_n10467,\t/a/ID_fun3 [1]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0101010000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2123|t/a/if_id/reg0_b0  (
    .a({_al_u2109_o,\t/a/if_id/n9 }),
    .b({\t/busarbitration/n3_placeOpt_3 ,\t/busarbitration/n3_placeOpt_3 }),
    .c({\t/busarbitration/instruction [12],\t/busarbitration/instruction [12]}),
    .clk(clock_pad),
    .d({i_data[12],i_data[12]}),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [12],open_n10481}),
    .q({open_n10485,\t/a/ID_fun3 [0]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u2124|_al_u596  (
    .a({\t/a/EX_fun7 [0],\t/a/ID_rs1$0$_placeOpt_12 }),
    .b({\t/a/EX_fun7 [1],\t/a/ID_rs1$1$_placeOpt_12 }),
    .c({\t/a/EX_fun7 [2],\t/a/regfile/regfile$4$ [27]}),
    .d({\t/a/EX_fun7 [3],\t/a/regfile/regfile$5$ [27]}),
    .f({_al_u2124_o,_al_u596_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(~0*D*C*B))"),
    //.LUTF1("~A*~B*C*D+A*~B*C*D"),
    //.LUTG0("(~A*~(~1*D*C*B))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0001010101010101),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b0101010101010101),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2125|_al_u2128  (
    .a({open_n10506,_al_u2126_o}),
    .b({\t/a/EX_fun7 [6],\t/a/EX_operation [2]}),
    .c({_al_u2124_o,\t/a/aluin/n35_lutinv }),
    .d({\t/a/EX_fun7 [5],\t/a/EX_fun3 [0]}),
    .e({\t/a/EX_fun7 [4],\t/a/EX_fun3 [1]}),
    .f({\t/a/aluin/n35_lutinv ,_al_u2128_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    //.LUTF1("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b0000000000110011),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b0011001100110011),
    .INIT_LUTG1(16'b0011001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2130|_al_u2406  (
    .a({\t/a/alu/n6 [31],open_n10529}),
    .b({_al_u2128_o,_al_u2128_o}),
    .d({open_n10534,\t/a/alu/n6 [17]}),
    .e({\t/a/EX_operation$0$_lutinv_placeOpt_2 ,\t/a/EX_operation$0$_lutinv_placeOpt_2 }),
    .f({_al_u2130_o,_al_u2406_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUTF1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0001000011110000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b0111000011110000),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2131|_al_u2436  (
    .a({\t/a/EX_A [14],\t/a/EX_A [15]}),
    .b({open_n10555,\t/a/EX_B [15]}),
    .c({open_n10556,\t/a/EX_operation [1]}),
    .d({\t/a/EX_A [15],\t/a/EX_operation [2]}),
    .e({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .f({\t/a/alu/n156_lutinv ,_al_u2436_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(A*~D))"),
    //.LUT1("(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111010),
    .INIT_LUT1(16'b1111101000001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2132|t/a/id_ex/reg7_b12  (
    .a({\t/a/EX_A [13],\t/a/EX_memstraddr [12]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel0_b12/B0 }),
    .clk(clock_pad),
    .d({\t/a/EX_A [12],_al_u1806_o}),
    .mi({open_n10592,\t/a/ID_memstraddr [12]}),
    .sr(rst_pad),
    .f({\t/a/alu/n158_lutinv ,\t/a/EX_A [12]}),
    .q({open_n10596,\t/a/EX_memstraddr [12]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    //.LUT1("~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .INIT_LUT0(16'b0001000111011101),
    .INIT_LUT1(16'b0001000111011101),
    .MODE("LOGIC"))
    \_al_u2133|_al_u2408  (
    .a({\t/a/alu/n156_lutinv ,\t/a/alu/n30_lutinv }),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n158_lutinv ,\t/a/alu/n28_lutinv }),
    .f({_al_u2133_o,_al_u2408_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~D*B*~C*~A+D*B*~C*~A+~D*B*C*~A+D*B*C*~A+~D*B*~C*A+D*B*~C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("D*~B*~C*~A+D*B*~C*~A+D*~B*C*~A+D*B*C*~A+D*~B*~C*A+D*B*~C*A+D*~B*C*A+D*B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111101011111010),
    .INIT_LUTF1(16'b1100110011001100),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b1111111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2134|t/a/id_ex/reg7_b10  (
    .a({open_n10619,\t/a/EX_memstraddr [10]}),
    .b({\t/a/EX_A [11],open_n10620}),
    .c({open_n10621,\t/a/aluin/sel0_b10/B0 }),
    .clk(clock_pad),
    .d({\t/a/EX_A [10],open_n10623}),
    .e({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u1806_o}),
    .mi({open_n10625,\t/a/ID_memstraddr [10]}),
    .sr(rst_pad),
    .f({\t/a/alu/n160_lutinv ,\t/a/EX_A [10]}),
    .q({open_n10640,\t/a/EX_memstraddr [10]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~A*B*~D+C*~A*B*~D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    //.LUTF1("A*D*~C*~B+A*D*C*~B+A*D*~C*B+A*D*C*B"),
    //.LUTG0("~C*A*B*~D+C*A*B*~D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    //.LUTG1("~A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+~A*D*C*~B+A*D*C*~B+~A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+~A*D*C*B+A*D*C*B"),
    .INIT_LUTF0(16'b1100110001000100),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b1100110010001000),
    .INIT_LUTG1(16'b1111111101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2135|_al_u2505  (
    .a({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o }),
    .b({open_n10641,_al_u2431_o}),
    .d({\t/a/EX_A [8],\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .e(\t/a/EX_A [9:8]),
    .f({\t/a/alu/n162_lutinv ,_al_u2505_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    //.LUT1("~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    .INIT_LUT0(16'b0101010100110011),
    .INIT_LUT1(16'b0010001001110111),
    .MODE("LOGIC"))
    \_al_u2136|_al_u2244  (
    .a({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/alu/n153_lutinv }),
    .b({\t/a/alu/n162_lutinv ,\t/a/alu/n151_lutinv }),
    .d({\t/a/alu/n160_lutinv ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2136_o,_al_u2244_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("~C*B*A*~D+C*B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG0("~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D"),
    //.LUTG1("~C*B*A*~D+C*B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*B*A*D+C*B*A*D"),
    .INIT_LUTF0(16'b1111111110101010),
    .INIT_LUTF1(16'b1101110110001000),
    .INIT_LUTG0(16'b0101010100000000),
    .INIT_LUTG1(16'b1101110110001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2137|_al_u2270  (
    .a({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .b({_al_u2136_o,open_n10688}),
    .d({_al_u2133_o,_al_u2269_o}),
    .e({open_n10693,\t/a/alu/n56_lutinv }),
    .f({_al_u2137_o,_al_u2270_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(A*~B))"),
    //.LUT1("(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001011110010),
    .INIT_LUT1(16'b1110111000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2138|t/a/id_ex/reg7_b7  (
    .a({\t/a/EX_A [7],\t/a/EX_memstraddr [7]}),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u1806_o}),
    .c({open_n10714,\t/a/aluin/sel0_b7/B0 }),
    .clk(clock_pad),
    .d({\t/a/EX_A [6],open_n10716}),
    .mi({open_n10727,\t/a/ID_memstraddr [7]}),
    .sr(rst_pad),
    .f({\t/a/alu/n164_lutinv ,\t/a/EX_A [7]}),
    .q({open_n10731,\t/a/EX_memstraddr [7]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~D*~C*~B+A*~D*C*~B+A*~D*~C*B+A*~D*C*B"),
    //.LUTF1("~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b0101010100000000),
    .INIT_LUTG0(16'b1111111111111111),
    .INIT_LUTG1(16'b1111111110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2139|t/a/id_ex/reg7_b4  (
    .a({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [4]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [5],_al_u1806_o}),
    .e({\t/a/EX_A [4],\t/a/aluin/sel0_b4/B0 }),
    .mi({open_n10738,\t/a/ID_memstraddr [4]}),
    .sr(rst_pad),
    .f({\t/a/alu/n166_lutinv ,\t/a/EX_A [4]}),
    .q({open_n10753,\t/a/EX_memstraddr [4]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    //.LUT1("~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)"),
    .INIT_LUT0(16'b1010111110100000),
    .INIT_LUT1(16'b0101010100001111),
    .MODE("LOGIC"))
    \_al_u2140|_al_u2260  (
    .a({\t/a/alu/n166_lutinv ,_al_u2140_o}),
    .c({\t/a/alu/n164_lutinv ,\t/a/EX_B [2]}),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,_al_u2136_o}),
    .f({_al_u2140_o,_al_u2260_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(A*~C))"),
    //.LUT1("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100001010),
    .INIT_LUT1(16'b1110010011100100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2141|t/a/id_ex/reg7_b3  (
    .a({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [3]}),
    .b({\t/a/EX_A [3],open_n10776}),
    .c({\t/a/EX_A [2],_al_u1806_o}),
    .clk(clock_pad),
    .d({open_n10778,\t/a/aluin/sel0_b3/B0 }),
    .mi({open_n10789,\t/a/ID_memstraddr [3]}),
    .sr(rst_pad),
    .f({\t/a/alu/n168_lutinv ,\t/a/EX_A [3]}),
    .q({open_n10793,\t/a/EX_memstraddr [3]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    //.LUT1("~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    .INIT_LUT0(16'b1010111110100000),
    .INIT_LUT1(16'b0001000110111011),
    .MODE("LOGIC"))
    \_al_u2143|_al_u2142  (
    .a({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [0]}),
    .b({\t/a/alu/n168_lutinv ,open_n10794}),
    .c({open_n10795,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n170_lutinv ,\t/a/EX_A [1]}),
    .f({_al_u2143_o,\t/a/alu/n170_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    //.LUT1("(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    .INIT_LUT0(16'b1110111001000100),
    .INIT_LUT1(16'b1111101000001010),
    .MODE("LOGIC"))
    \_al_u2144|_al_u2384  (
    .a({_al_u2140_o,\t/a/EX_B [2]}),
    .b({open_n10816,_al_u2383_o}),
    .c({\t/a/EX_B [2],open_n10817}),
    .d({_al_u2143_o,_al_u2332_o}),
    .f({_al_u2144_o,_al_u2384_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0011000000110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2146|_al_u2161  (
    .b({open_n10840,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_operation$0$_lutinv_placeOpt_2 ,\t/a/EX_operation$0$_lutinv_placeOpt_2 }),
    .d({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,open_n10843}),
    .f({_al_u2146_o,_al_u2161_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~B)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~B)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0011000000110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0011000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2147|_al_u2313  (
    .b({_al_u2145_o,open_n10864}),
    .c({_al_u2146_o,_al_u2146_o}),
    .d({open_n10867,_al_u2312_o}),
    .f({_al_u2147_o,_al_u2313_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(A*~D))"),
    //.LUT1("(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011111010),
    .INIT_LUT1(16'b1011101110001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2148|t/a/id_ex/reg7_b22  (
    .a({\t/a/EX_A [22],\t/a/EX_memstraddr [22]}),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,open_n10890}),
    .c({open_n10891,\t/a/aluin/sel0_b22/B0 }),
    .clk(clock_pad),
    .d({\t/a/EX_A [23],_al_u1806_o}),
    .mi({open_n10903,\t/a/ID_memstraddr [22]}),
    .sr(rst_pad),
    .f({\t/a/alu/n148_lutinv ,\t/a/EX_A [22]}),
    .q({open_n10907,\t/a/EX_memstraddr [22]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(A*~B))"),
    //.LUT1("(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100100010),
    .INIT_LUT1(16'b1110111000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2149|t/a/id_ex/reg7_b21  (
    .a({\t/a/EX_A [21],\t/a/EX_memstraddr [21]}),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u1806_o}),
    .clk(clock_pad),
    .d({\t/a/EX_A [20],\t/a/aluin/sel0_b21/B0 }),
    .mi({open_n10921,\t/a/ID_memstraddr [21]}),
    .sr(rst_pad),
    .f({\t/a/alu/n150_lutinv ,\t/a/EX_A [21]}),
    .q({open_n10925,\t/a/EX_memstraddr [21]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D"),
    .INIT_LUTF0(16'b0101000001011111),
    .INIT_LUTF1(16'b1111000011111111),
    .INIT_LUTG0(16'b0101000001011111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2150|_al_u2237  (
    .a({open_n10926,\t/a/alu/n161_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n148_lutinv ,\t/a/alu/n159_lutinv }),
    .e({\t/a/alu/n150_lutinv ,open_n10931}),
    .f({_al_u2150_o,_al_u2237_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~C*~B*~D+A*~C*B*~D+A*~C*~B*D+A*~C*B*D"),
    //.LUTF1("(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)"),
    //.LUTG0("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG1("(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000001010),
    .INIT_LUTF1(16'b1011101110001000),
    .INIT_LUTG0(16'b1111111111111111),
    .INIT_LUTG1(16'b1011101110001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2151|t/a/id_ex/reg7_b19  (
    .a({\t/a/EX_A [18],\t/a/EX_memstraddr [19]}),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,open_n10952}),
    .c({open_n10953,_al_u1806_o}),
    .clk(clock_pad),
    .d({\t/a/EX_A [19],open_n10955}),
    .e({open_n10956,\t/a/aluin/sel0_b19/B0 }),
    .mi({open_n10958,\t/a/ID_memstraddr [19]}),
    .sr(rst_pad),
    .f({\t/a/alu/n152_lutinv ,\t/a/EX_A [19]}),
    .q({open_n10973,\t/a/EX_memstraddr [19]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(A*~B))"),
    //.LUT1("(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100100010),
    .INIT_LUT1(16'b1010101011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2152|t/a/id_ex/reg7_b17  (
    .a({\t/a/EX_A [16],\t/a/EX_memstraddr [17]}),
    .b({\t/a/EX_A [17],_al_u1806_o}),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel0_b17/B0 }),
    .mi({open_n10987,\t/a/ID_memstraddr [17]}),
    .sr(rst_pad),
    .f({\t/a/alu/n154_lutinv ,\t/a/EX_A [17]}),
    .q({open_n10991,\t/a/EX_memstraddr [17]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    //.LUT1("~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    .INIT_LUT0(16'b0010001001110111),
    .INIT_LUT1(16'b0001000110111011),
    .MODE("LOGIC"))
    \_al_u2153|_al_u2221  (
    .a({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .b({\t/a/alu/n152_lutinv ,\t/a/alu/n152_lutinv }),
    .d({\t/a/alu/n154_lutinv ,\t/a/alu/n150_lutinv }),
    .f({_al_u2153_o,_al_u2221_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    //.LUT1("(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)"),
    .INIT_LUT0(16'b1010110010101100),
    .INIT_LUT1(16'b1011101110001000),
    .MODE("LOGIC"))
    \_al_u2154|_al_u2265  (
    .a({_al_u2153_o,_al_u2133_o}),
    .b({\t/a/EX_B [2],_al_u2153_o}),
    .c({open_n11014,\t/a/EX_B [2]}),
    .d({_al_u2150_o,open_n11017}),
    .f({_al_u2154_o,_al_u2265_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*~(A*~D))"),
    //.LUTF1("~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~(~C*~(A*~D))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011111010),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000011111010),
    .INIT_LUTG1(16'b1111111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2155|t/a/id_ex/reg7_b27  (
    .a({open_n11036,\t/a/EX_memstraddr [27]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel0_b27/B0 }),
    .clk(clock_pad),
    .d({\t/a/EX_A [26],_al_u1806_o}),
    .e({\t/a/EX_A [27],open_n11040}),
    .mi({open_n11042,\t/a/ID_memstraddr [27]}),
    .sr(rst_pad),
    .f({\t/a/alu/n144_lutinv ,\t/a/EX_A [27]}),
    .q({open_n11057,\t/a/EX_memstraddr [27]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1011100010111000),
    .MODE("LOGIC"))
    \_al_u2156|_al_u649  (
    .a({\t/a/EX_A [24],\t/a/ID_rs1$0$_placeOpt_15 }),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/ID_rs1$1$_placeOpt_15 }),
    .c({\t/a/EX_A [25],\t/a/regfile/regfile$4$ [24]}),
    .d({open_n11060,\t/a/regfile/regfile$5$ [24]}),
    .f({\t/a/alu/n146_lutinv ,_al_u649_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+~A*C*B*D"),
    //.LUTF1("~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)"),
    //.LUTG0("~A*~C*B*~D+~A*C*B*~D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG1("~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)"),
    .INIT_LUTF0(16'b0111011101110111),
    .INIT_LUTF1(16'b0011001101010101),
    .INIT_LUTG0(16'b0100010001000100),
    .INIT_LUTG1(16'b0011001101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2157|_al_u2224  (
    .a({\t/a/alu/n144_lutinv ,\t/a/alu/n148_lutinv }),
    .b({\t/a/alu/n146_lutinv ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n11083}),
    .e({open_n11084,\t/a/alu/n146_lutinv }),
    .f({_al_u2157_o,_al_u2224_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(A*~C))"),
    //.LUTF1("D*~B*C*~A+D*B*C*~A+D*~B*C*A+D*B*C*A"),
    //.LUTG0("~(~D*~(A*~C))"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+D*~B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+D*~B*C*A+D*B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100001010),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111111100001010),
    .INIT_LUTG1(16'b1111111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2158|t/a/id_ex/reg7_b28  (
    .a({open_n11105,\t/a/EX_memstraddr [28]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u1806_o}),
    .clk(clock_pad),
    .d({\t/a/EX_A [28],\t/a/aluin/sel0_b28/B0 }),
    .e({\t/a/EX_A [29],open_n11109}),
    .mi({open_n11111,\t/a/ID_memstraddr [28]}),
    .sr(rst_pad),
    .f({\t/a/alu/n142_lutinv ,\t/a/EX_A [28]}),
    .q({open_n11126,\t/a/EX_memstraddr [28]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("(~1*~(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)))"),
    .INIT_LUT0(16'b1111001111110101),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2159 (
    .a({\t/a/EX_A [30],\t/a/EX_A [31]}),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [30]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_A [31],\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .mi({open_n11139,\t/a/EX_B [2]}),
    .fx({open_n11144,_al_u2159_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~(D*B)*C)*~(0*A))"),
    //.LUT1("(~(~(B*D)*C)*~(1*A))"),
    .INIT_LUT0(16'b1100111100001111),
    .INIT_LUT1(16'b0100010100000101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2160 (
    .a({_al_u2157_o,_al_u2157_o}),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/alu/n142_lutinv }),
    .c({_al_u2159_o,_al_u2159_o}),
    .d({\t/a/alu/n142_lutinv ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .mi({open_n11159,\t/a/EX_B [2]}),
    .fx({open_n11164,\t/a/alu/n204_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~A*C*~B+D*~A*C*~B+~D*A*C*~B+D*A*C*~B+~D*~A*C*B+D*~A*C*B"),
    //.LUTF1("~D*B*C*~A+D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("~D*~A*C*B+D*~A*C*B"),
    //.LUTG1("~D*B*C*~A+D*B*C*~A"),
    .INIT_LUTF0(16'b0111000001110000),
    .INIT_LUTF1(16'b1110000011100000),
    .INIT_LUTG0(16'b0100000001000000),
    .INIT_LUTG1(16'b0100000001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2162|_al_u2328  (
    .a({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 ,_al_u2137_o}),
    .b({\t/a/alu/n204_lutinv ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }),
    .c({_al_u2161_o,_al_u2161_o}),
    .e({_al_u2154_o,_al_u2154_o}),
    .f({_al_u2162_o,_al_u2328_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2163 (
    .a({\t/a/alu/n5 [31],\t/a/alu/n5 [31]}),
    .b({_al_u2147_o,_al_u2147_o}),
    .c({_al_u2162_o,_al_u2162_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n11203,\t/a/EX_operation$0$_lutinv_placeOpt_2 }),
    .fx({open_n11208,_al_u2163_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~C*~(A*~B))"),
    //.LUT1("(~A*~D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001011110010),
    .INIT_LUT1(16'b0000000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2164|t/a/id_ex/reg7_b31  (
    .a({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [31]}),
    .b({open_n11211,_al_u1806_o}),
    .c({\t/a/EX_A [31],\t/a/aluin/sel0_b31/B0 }),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n11213}),
    .mi({open_n11224,\t/a/ID_memstraddr [31]}),
    .sr(rst_pad),
    .f({\t/a/alu/n56_lutinv ,\t/a/EX_A [31]}),
    .q({open_n11228,\t/a/EX_memstraddr [31]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~D*C*A))"),
    //.LUTF1("(~D*~A)"),
    //.LUTG0("(B*~(~1*~D*C*A))"),
    //.LUTG1("(~D*~A)"),
    .INIT_LUTF0(16'b1100110001001100),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2168|_al_u2166  (
    .a({_al_u2166_o,\t/a/alu/n56_lutinv }),
    .b({open_n11229,_al_u2165_o}),
    .c({open_n11230,_al_u2161_o}),
    .d({\t/a/EX_operation [1],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .e({open_n11233,\t/a/EX_B [2]}),
    .f({_al_u2168_o,_al_u2166_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(B*(D*~(A)*~(C)+~(D)*A*~(C)+D*A*~(C)+D*A*C))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b1000110000001000),
    .MODE("LOGIC"))
    \_al_u2170|_al_u2165  (
    .a({\t/a/EX_B [31],\t/a/EX_A [31]}),
    .b({_al_u2169_o,\t/a/EX_B [31]}),
    .c({\t/a/EX_operation$0$_lutinv_placeOpt_1 ,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .d({\t/a/EX_A [31],\t/a/EX_operation [2]}),
    .f({_al_u2170_o,_al_u2165_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("(~C*~(~A*D))"),
    //.LUTG0("0"),
    //.LUTG1("(~C*~(~A*D))"),
    .INIT_LUTF0(16'b1111111101010101),
    .INIT_LUTF1(16'b0000101000001111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000101000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2172|_al_u2369  (
    .a({\t/a/EX_operation$0$_lutinv_placeOpt_5 ,\t/a/alu/n6 [20]}),
    .c({_al_u2128_o,open_n11276}),
    .d({\t/a/alu/n6 [30],\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .e({open_n11279,_al_u2128_o}),
    .f({_al_u2172_o,_al_u2369_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~D*(B@A)))"),
    //.LUT1("(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .INIT_LUT0(16'b1111000010010000),
    .INIT_LUT1(16'b1110111000100010),
    .MODE("LOGIC"))
    \_al_u2173|_al_u2455  (
    .a(\t/a/EX_A [14:13]),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [13]}),
    .c({open_n11300,_al_u2431_o}),
    .d({\t/a/EX_A [13],\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .f({\t/a/alu/n157_lutinv ,_al_u2455_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    //.LUT1("~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .INIT_LUT0(16'b1010111110100000),
    .INIT_LUT1(16'b0001000111011101),
    .MODE("LOGIC"))
    \_al_u2175|_al_u2174  (
    .a({\t/a/alu/n157_lutinv ,\t/a/EX_A [11]}),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n11321}),
    .c({open_n11322,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n159_lutinv ,\t/a/EX_A [12]}),
    .f({_al_u2175_o,\t/a/alu/n159_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~D*(B@A)))"),
    //.LUT1("(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    .INIT_LUT0(16'b1111000010010000),
    .INIT_LUT1(16'b1111101000001010),
    .MODE("LOGIC"))
    \_al_u2176|_al_u2485  (
    .a({\t/a/EX_A [10],\t/a/EX_A [10]}),
    .b({open_n11343,\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2431_o}),
    .d({\t/a/EX_A [9],\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .f({\t/a/alu/n161_lutinv ,_al_u2485_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b1101110110001000),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b1101110110001000),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2178|_al_u2177  (
    .a({\t/a/alu/n163_lutinv ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .b({open_n11364,\t/a/EX_A [7]}),
    .d({\t/a/alu/n161_lutinv ,\t/a/EX_A [8]}),
    .e({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n11369}),
    .f({_al_u2178_o,\t/a/alu/n163_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+D*C*~B*A"),
    //.LUTF1("~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    //.LUTG0("~D*~C*B*~A+D*~C*B*~A+~D*C*B*~A+D*C*B*~A+~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+D*C*~B*A+~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    //.LUTG1("~D*~C*~B*~A+D*~C*~B*~A+~D*C*~B*~A+D*C*~B*~A+~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+D*C*~B*A+~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    .INIT_LUTF0(16'b0010001000100010),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1011101110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2179|_al_u2282  (
    .a({_al_u2178_o,_al_u2194_o}),
    .b({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .e({_al_u2175_o,_al_u2175_o}),
    .f({_al_u2179_o,_al_u2282_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~C*~B*~D+A*~C*B*~D+A*~C*~B*D+A*~C*B*D"),
    //.LUTF1("A*~D*~C*B+A*D*~C*B+A*~D*C*B+A*D*C*B"),
    //.LUTG0("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG1("~A*~D*~C*~B+~A*D*~C*~B+~A*~D*C*~B+~A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000001010),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1111111111111111),
    .INIT_LUTG1(16'b1101110111011101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2180|t/a/id_ex/reg7_b6  (
    .a({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [6]}),
    .b({\t/a/EX_A [5],open_n11416}),
    .c({open_n11417,_al_u1806_o}),
    .clk(clock_pad),
    .e({\t/a/EX_A [6],\t/a/aluin/sel0_b6/B0 }),
    .mi({open_n11422,\t/a/ID_memstraddr [6]}),
    .sr(rst_pad),
    .f({\t/a/alu/n165_lutinv ,\t/a/EX_A [6]}),
    .q({open_n11437,\t/a/EX_memstraddr [6]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D"),
    //.LUTF1("~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("A*~C*~B*~D+A*C*~B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0011001100010001),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0011001100100010),
    .INIT_LUTG1(16'b1111111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2181|_al_u2546  (
    .a({open_n11438,\t/a/EX_A [4]}),
    .b({open_n11439,\t/a/EX_operation [1]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,open_n11440}),
    .d({\t/a/EX_A [3],\t/a/EX_operation [0]}),
    .e({\t/a/EX_A [4],\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .f({\t/a/alu/n167_lutinv ,_al_u2546_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D"),
    .INIT_LUTF0(16'b1111111100000000),
    .INIT_LUTF1(16'b1111000011111111),
    .INIT_LUTG0(16'b1010101010101010),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2182|_al_u2277  (
    .a({open_n11463,_al_u2182_o}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n11466}),
    .d({\t/a/alu/n165_lutinv ,_al_u2178_o}),
    .e({\t/a/alu/n167_lutinv ,\t/a/EX_B [2]}),
    .f({_al_u2182_o,_al_u2277_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~A*D*~C*~B+A*D*~C*~B+~A*D*C*~B+A*D*C*~B+~A*D*~C*B+A*D*~C*B+~A*D*C*B+A*D*C*B"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("A*~D*~C*~B+A*D*~C*~B+A*~D*C*~B+A*D*C*~B+A*~D*~C*B+A*D*~C*B+A*~D*C*B+A*D*C*B"),
    .INIT_LUTF0(16'b0101000001010000),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b1111101011111010),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2183|_al_u2559  (
    .a({\t/a/EX_A [1],\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .c({open_n11491,\t/a/EX_A [2]}),
    .d({\t/a/EX_A [2],open_n11494}),
    .e({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [3]}),
    .f({\t/a/alu/n169_lutinv ,\t/a/alu/n45_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    //.LUT1("(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)"),
    .INIT_LUT0(16'b0101010100110011),
    .INIT_LUT1(16'b1011101110001000),
    .MODE("LOGIC"))
    \_al_u2186|_al_u2185  (
    .a({_al_u2185_o,_al_u2184_o}),
    .b({\t/a/EX_B [2],\t/a/alu/n169_lutinv }),
    .d({_al_u2182_o,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2186_o,_al_u2185_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~A*~(~0*B))"),
    //.LUTF1("(B*~A)"),
    //.LUTG0("(D*~C*~A*~(~1*B))"),
    //.LUTG1("(B*~A)"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b0000010100000000),
    .INIT_LUTG1(16'b0100010001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2188|_al_u2203  (
    .a({_al_u2187_o,_al_u2188_o}),
    .b({_al_u2146_o,\t/a/alu/n5 [30]}),
    .c({open_n11537,_al_u2202_o}),
    .d({open_n11540,_al_u2128_o}),
    .e({open_n11541,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .f({_al_u2188_o,_al_u2203_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~C*B*~D+A*C*B*~D"),
    //.LUTF1("D*~B*C*~A+D*B*C*~A+D*~B*C*A+D*B*C*A"),
    //.LUTG0("~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+A*~C*B*D+A*C*B*D"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+D*~B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+D*~B*C*A+D*B*C*A"),
    .INIT_LUTF0(16'b0000000010001000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1000100011001100),
    .INIT_LUTG1(16'b1111111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2189|_al_u2363  (
    .a({open_n11562,\t/a/EX_A [21]}),
    .b({open_n11563,_al_u2169_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,open_n11564}),
    .d({\t/a/EX_A [21],\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .e({\t/a/EX_A [22],\t/a/EX_B [21]}),
    .f({\t/a/alu/n149_lutinv ,_al_u2363_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*C*~D+A*B*C*~D"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000000011000000),
    .INIT_LUTF1(16'b0000000010101010),
    .INIT_LUTG0(16'b1100000011110000),
    .INIT_LUTG1(16'b1111111110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2190|_al_u2388  (
    .a({\t/a/EX_A [20],open_n11587}),
    .b({open_n11588,\t/a/EX_B [19]}),
    .c({open_n11589,_al_u2169_o}),
    .d({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .e({\t/a/EX_A [19],\t/a/EX_A [19]}),
    .f({\t/a/alu/n151_lutinv ,_al_u2388_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    //.LUT1("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT_LUT0(16'b0011010100110101),
    .INIT_LUT1(16'b0101001101010011),
    .MODE("LOGIC"))
    \_al_u2191|_al_u2247  (
    .a({\t/a/alu/n151_lutinv ,\t/a/alu/n147_lutinv }),
    .b({\t/a/alu/n149_lutinv ,\t/a/alu/n149_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2191_o,_al_u2247_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D"),
    //.LUTG0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111110101010),
    .INIT_LUTF1(16'b0000000010101010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1111111110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2192|t/a/id_ex/reg7_b18  (
    .a({\t/a/EX_A [18],\t/a/EX_memstraddr [18]}),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel0_b18/B0 }),
    .e({\t/a/EX_A [17],_al_u1806_o}),
    .mi({open_n11640,\t/a/ID_memstraddr [18]}),
    .sr(rst_pad),
    .f({\t/a/alu/n153_lutinv ,\t/a/EX_A [18]}),
    .q({open_n11655,\t/a/EX_memstraddr [18]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2193|_al_u2425  (
    .a({open_n11656,\t/a/EX_A [16]}),
    .b({\t/a/EX_A [15],\t/a/EX_B [16]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [16],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n155_lutinv ,_al_u2425_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    //.LUT1("~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .INIT_LUT0(16'b1100101011001010),
    .INIT_LUT1(16'b0001000111011101),
    .MODE("LOGIC"))
    \_al_u2194|_al_u2195  (
    .a({\t/a/alu/n153_lutinv ,_al_u2191_o}),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,_al_u2194_o}),
    .c({open_n11677,\t/a/EX_B [2]}),
    .d({\t/a/alu/n155_lutinv ,open_n11680}),
    .f({_al_u2194_o,_al_u2195_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1011101110001000),
    .MODE("LOGIC"))
    \_al_u2196|_al_u2308  (
    .a({\t/a/EX_A [25],\t/a/EX_A [25]}),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [25]}),
    .c({open_n11699,_al_u2169_o}),
    .d({\t/a/EX_A [26],\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .f({\t/a/alu/n145_lutinv ,_al_u2308_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*C*~D+A*B*C*~D"),
    //.LUTF1("~A*C*~D*~B+A*C*~D*~B+~A*C*~D*B+A*C*~D*B"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*C*~D*~B+A*C*~D*~B+~A*~C*D*~B+A*~C*D*~B+~A*C*D*~B+A*C*D*~B+~A*C*~D*B+A*C*~D*B+~A*~C*D*B+A*~C*D*B+~A*C*D*B+A*C*D*B"),
    .INIT_LUTF0(16'b0000000011000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1100000011110000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2197|_al_u2337  (
    .b({open_n11722,\t/a/EX_B [23]}),
    .c({\t/a/EX_A [24],_al_u2169_o}),
    .d({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .e({\t/a/EX_A [23],\t/a/EX_A [23]}),
    .f({\t/a/alu/n147_lutinv ,_al_u2337_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)"),
    //.LUT1("~(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)"),
    .INIT_LUT0(16'b0100010001110111),
    .INIT_LUT1(16'b0100010001110111),
    .MODE("LOGIC"))
    \_al_u2198|_al_u2216  (
    .a({\t/a/alu/n147_lutinv ,\t/a/alu/n168_lutinv }),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n145_lutinv ,\t/a/alu/n166_lutinv }),
    .f({_al_u2198_o,_al_u2216_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*B*D*~A+C*B*D*~A"),
    //.LUTF1("~A*B*C*~D+A*B*C*~D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~C*~B*D*~A+C*~B*D*~A+~C*B*D*~A+C*B*D*~A+~C*B*D*A+C*B*D*A"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0100010000000000),
    .INIT_LUTF1(16'b1100000011000000),
    .INIT_LUTG0(16'b1101110100000000),
    .INIT_LUTG1(16'b1100111111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2199|_al_u2274  (
    .a({open_n11767,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .b({\t/a/EX_A [27],\t/a/EX_B [27]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,open_n11768}),
    .d({open_n11771,_al_u2169_o}),
    .e(\t/a/EX_A [28:27]),
    .f({\t/a/alu/n143_lutinv ,_al_u2274_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("((B*~(C)*~(0)+B*C*~(0)+~(B)*C*0+B*C*0)*~(A)*~(D)+(B*~(C)*~(0)+B*C*~(0)+~(B)*C*0+B*C*0)*A*~(D)+~((B*~(C)*~(0)+B*C*~(0)+~(B)*C*0+B*C*0))*A*D+(B*~(C)*~(0)+B*C*~(0)+~(B)*C*0+B*C*0)*A*D)"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*B*~C*D+A*B*C*D"),
    //.LUTG0("((B*~(C)*~(1)+B*C*~(1)+~(B)*C*1+B*C*1)*~(A)*~(D)+(B*~(C)*~(1)+B*C*~(1)+~(B)*C*1+B*C*1)*A*~(D)+~((B*~(C)*~(1)+B*C*~(1)+~(B)*C*1+B*C*1))*A*D+(B*~(C)*~(1)+B*C*~(1)+~(B)*C*1+B*C*1)*A*D)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1010101011001100),
    .INIT_LUTF1(16'b1000100011011101),
    .INIT_LUTG0(16'b1010101011110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2201|_al_u2200  (
    .a({\t/a/EX_B [2],\t/a/alu/n143_lutinv }),
    .b({_al_u2198_o,\t/a/EX_A [30]}),
    .c({open_n11792,\t/a/EX_A [29]}),
    .d({\t/a/alu/n173_lutinv ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2201_o,\t/a/alu/n173_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(C*~B*~(D*A))"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0001000000110000),
    .MODE("LOGIC"))
    \_al_u2202|_al_u2341  (
    .a({_al_u2195_o,_al_u2195_o}),
    .b({_al_u2201_o,_al_u2179_o}),
    .c({_al_u2161_o,_al_u2161_o}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }),
    .f({_al_u2202_o,_al_u2341_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~D*A*B+C*~D*A*B+~C*D*A*B+C*D*A*B"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("~C*~D*~A*~B+C*~D*~A*~B+~C*D*~A*~B+C*D*~A*~B+~C*~D*~A*B+C*~D*~A*B+~C*D*~A*B+C*D*~A*B+~C*~D*A*B+C*~D*A*B+~C*D*A*B+C*D*A*B"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b1010101010101010),
    .INIT_LUTG0(16'b1101110111011101),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2205|_al_u2204  (
    .a({\t/a/alu/n17_lutinv ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .b({open_n11835,\t/a/EX_A [31]}),
    .e({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [30]}),
    .f({\t/a/alu/n57_lutinv ,\t/a/alu/n17_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D)*~(B)+~A*D*~(B)+~(~A)*D*B+~A*D*B)"),
    //.LUT1("(~A*D)"),
    .INIT_LUT0(16'b0010001011101110),
    .INIT_LUT1(16'b0101010100000000),
    .MODE("LOGIC"))
    \_al_u2206|_al_u2287  (
    .a({\t/a/EX_B [2],_al_u2286_o}),
    .b({open_n11862,\t/a/EX_B [2]}),
    .d({\t/a/alu/n57_lutinv ,\t/a/alu/n57_lutinv }),
    .f({\t/a/alu/n106_lutinv ,_al_u2287_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D"),
    //.LUTF1("(~C*B)"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTG1("(~C*B)"),
    .INIT_LUTF0(16'b0011000000110000),
    .INIT_LUTF1(16'b0000110000001100),
    .INIT_LUTG0(16'b0011111100111111),
    .INIT_LUTG1(16'b0000110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2207|_al_u2347  (
    .b({\t/a/alu/n106_lutinv ,\t/a/alu/n106_lutinv }),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }),
    .e({open_n11891,_al_u2346_o}),
    .f({\t/a/alu/n138_lutinv ,_al_u2347_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*~A*C+D*~B*~A*C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    //.LUTG0("~D*B*~A*C+D*B*~A*C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b1110000011100000),
    .INIT_LUTG1(16'b0010001000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2209|_al_u2208  (
    .a({\t/a/alu/n138_lutinv ,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .b({\t/a/EX_operation [1],\t/a/EX_B [30]}),
    .c({open_n11912,\t/a/EX_operation [2]}),
    .d({_al_u2208_o,open_n11915}),
    .e({_al_u2161_o,\t/a/EX_A [30]}),
    .f({_al_u2209_o,_al_u2208_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(B*(D*~(A)*~(C)+~(D)*A*~(C)+D*A*~(C)+D*A*C))"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1000110000001000),
    .MODE("LOGIC"))
    \_al_u2210|_al_u2234  (
    .a({\t/a/EX_B [30],\t/a/EX_A [29]}),
    .b({_al_u2169_o,\t/a/EX_B [29]}),
    .c({\t/a/EX_operation$0$_lutinv_placeOpt_4 ,_al_u2169_o}),
    .d({\t/a/EX_A [30],\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .f({_al_u2210_o,_al_u2234_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~D*A))"),
    //.LUT1("(~B*~(~D*A))"),
    .INIT_LUT0(16'b0011001100010001),
    .INIT_LUT1(16'b0011001100010001),
    .MODE("LOGIC"))
    \_al_u2212|_al_u2356  (
    .a({\t/a/alu/n6 [29],\t/a/alu/n6 [21]}),
    .b({_al_u2128_o,_al_u2128_o}),
    .d({\t/a/EX_operation$0$_lutinv_placeOpt_4 ,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .f({_al_u2212_o,_al_u2356_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D"),
    //.LUTG1("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b1111000011111111),
    .INIT_LUTF1(16'b0101111101011111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0101000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2213|_al_u2214  (
    .a({\t/a/alu/n160_lutinv ,open_n11978}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({open_n11983,\t/a/alu/n162_lutinv }),
    .e({\t/a/alu/n158_lutinv ,\t/a/alu/n164_lutinv }),
    .f({_al_u2213_o,_al_u2214_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1100110011001100),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2215|_al_u2299  (
    .b({_al_u2213_o,open_n12006}),
    .c({open_n12007,\t/a/EX_B [2]}),
    .d({_al_u2214_o,_al_u2222_o}),
    .e({\t/a/EX_B [2],_al_u2213_o}),
    .f({_al_u2215_o,_al_u2299_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    //.LUT1("~(~A*~(D)*~(C)+~A*D*~(C)+~(~A)*D*C+~A*D*C)"),
    .INIT_LUT0(16'b1101110110001000),
    .INIT_LUT1(16'b0000101011111010),
    .MODE("LOGIC"))
    \_al_u2218|_al_u2294  (
    .a({_al_u2216_o,\t/a/EX_B [2]}),
    .b({open_n12030,_al_u2216_o}),
    .c({\t/a/EX_B [2],open_n12031}),
    .d({\t/a/alu/n202_lutinv ,_al_u2214_o}),
    .f({_al_u2218_o,_al_u2294_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~C*~D*~(~0*A))"),
    //.LUTF1("(A*~B)"),
    //.LUTG0("(B*~C*~D*~(~1*A))"),
    //.LUTG1("(A*~B)"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b0010001000100010),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0010001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2220|_al_u2227  (
    .a({_al_u2146_o,\t/a/alu/n5 [29]}),
    .b({_al_u2219_o,_al_u2128_o}),
    .c({open_n12052,_al_u2226_o}),
    .d({open_n12055,_al_u2220_o}),
    .e({open_n12056,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .f({_al_u2220_o,_al_u2227_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    //.LUT1("~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    .INIT_LUT0(16'b1101110110001000),
    .INIT_LUT1(16'b0101000001011111),
    .MODE("LOGIC"))
    \_al_u2222|_al_u2223  (
    .a({\t/a/alu/n156_lutinv ,\t/a/EX_B [2]}),
    .b({open_n12077,_al_u2222_o}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n12078}),
    .d({\t/a/alu/n154_lutinv ,_al_u2221_o}),
    .f({_al_u2222_o,_al_u2223_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(0)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(0)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*0+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*0)"),
    //.LUT1("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(1)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(1)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*1+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*1)"),
    .INIT_LUT0(16'b0011001100001111),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2225 (
    .a({_al_u2224_o,_al_u2224_o}),
    .b({\t/a/alu/n144_lutinv ,\t/a/alu/n144_lutinv }),
    .c({\t/a/alu/n142_lutinv ,\t/a/alu/n142_lutinv }),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .mi({open_n12111,\t/a/EX_B [2]}),
    .fx({open_n12116,_al_u2225_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~A*C*~B+D*~A*C*~B+~D*A*C*~B+D*A*C*~B+~D*~A*C*B+D*~A*C*B"),
    //.LUTF1("~D*~B*A*~C+D*~B*A*~C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTG0("~D*~A*C*B+D*~A*C*B"),
    //.LUTG1("~D*~B*A*~C+D*~B*A*~C"),
    .INIT_LUTF0(16'b0111000001110000),
    .INIT_LUTF1(16'b1010001010100010),
    .INIT_LUTG0(16'b0100000001000000),
    .INIT_LUTG1(16'b0000001000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2226|_al_u2354  (
    .a({_al_u2161_o,_al_u2215_o}),
    .b({_al_u2225_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 }),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 ,_al_u2161_o}),
    .e({_al_u2223_o,_al_u2223_o}),
    .f({_al_u2226_o,_al_u2354_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~((~D*B))*~(C)+A*(~D*B)*~(C)+~(A)*(~D*B)*C+A*(~D*B)*C)"),
    //.LUT1("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT_LUT0(16'b1111010100110101),
    .INIT_LUT1(16'b1110001011100010),
    .MODE("LOGIC"))
    \_al_u2228|_al_u2229  (
    .a({\t/a/EX_A [29],\t/a/alu/n18_lutinv }),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [31]}),
    .c({\t/a/EX_A [30],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({open_n12145,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({\t/a/alu/n18_lutinv ,_al_u2229_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("(~C*A)"),
    //.LUTG0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTG1("(~C*A)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2231|_al_u2360  (
    .a({\t/a/alu/n105_lutinv ,open_n12164}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 }),
    .d({open_n12169,_al_u2359_o}),
    .e({open_n12170,\t/a/alu/n105_lutinv }),
    .f({\t/a/alu/n137_lutinv ,_al_u2360_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*~A*C+D*~B*~A*C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTF1("~A*~D*~C*~B+~A*D*~C*~B+~A*~D*C*~B+~A*D*C*~B"),
    //.LUTG0("~D*B*~A*C+D*B*~A*C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTG1("~A*~D*~C*~B+~A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b1110000011100000),
    .INIT_LUTG1(16'b0011000100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2233|_al_u2232  (
    .a({_al_u2232_o,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .b({\t/a/EX_operation [1],\t/a/EX_B [29]}),
    .c({_al_u2161_o,\t/a/EX_operation [2]}),
    .e({\t/a/alu/n137_lutinv ,\t/a/EX_A [29]}),
    .f({_al_u2233_o,_al_u2232_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~C*D))"),
    //.LUT1("(~A*~(~C*D))"),
    .INIT_LUT0(16'b0101000001010101),
    .INIT_LUT1(16'b0101000001010101),
    .MODE("LOGIC"))
    \_al_u2236|_al_u2343  (
    .a({_al_u2128_o,_al_u2128_o}),
    .c({\t/a/EX_operation$0$_lutinv_placeOpt_4 ,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .d({\t/a/alu/n6 [28],\t/a/alu/n6 [22]}),
    .f({_al_u2236_o,_al_u2343_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*~C*D+A*B*~C*D"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D"),
    .INIT_LUTF0(16'b0000101000001010),
    .INIT_LUTF1(16'b0011001111111111),
    .INIT_LUTG0(16'b1111101011111010),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2238|_al_u2239  (
    .a({open_n12237,_al_u2237_o}),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n12238}),
    .c({open_n12239,\t/a/EX_B [2]}),
    .d({\t/a/alu/n165_lutinv ,open_n12242}),
    .e({\t/a/alu/n163_lutinv ,_al_u2238_o}),
    .f({_al_u2238_o,_al_u2239_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b1111010100000000),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b1111010111111111),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2240|_al_u2241  (
    .a({\t/a/alu/n169_lutinv ,_al_u2184_o}),
    .c({open_n12265,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n167_lutinv ,\t/a/EX_B [2]}),
    .e({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,_al_u2240_o}),
    .f({_al_u2240_o,_al_u2241_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b1110111001000100),
    .MODE("LOGIC"))
    \_al_u2242|_al_u2367  (
    .a({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,_al_u2246_o}),
    .b({_al_u2239_o,_al_u2239_o}),
    .c({open_n12288,_al_u2161_o}),
    .d({_al_u2241_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2242_o,_al_u2367_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~D)"),
    //.LUT1("(B*~C)"),
    .INIT_LUT0(16'b0000000011001100),
    .INIT_LUT1(16'b0000110000001100),
    .MODE("LOGIC"))
    \_al_u2243|_al_u2263  (
    .b({_al_u2146_o,_al_u2146_o}),
    .c({_al_u2242_o,open_n12311}),
    .d({open_n12314,_al_u2262_o}),
    .f({_al_u2243_o,_al_u2263_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A"),
    .INIT_LUTF0(16'b1010101011001100),
    .INIT_LUTF1(16'b1111010111110101),
    .INIT_LUTG0(16'b1010101011001100),
    .INIT_LUTG1(16'b0000010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2245|_al_u2246  (
    .a({\t/a/alu/n155_lutinv ,_al_u2245_o}),
    .b({open_n12333,_al_u2244_o}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n12334}),
    .d({open_n12337,\t/a/EX_B [2]}),
    .e({\t/a/alu/n157_lutinv ,open_n12338}),
    .f({_al_u2245_o,_al_u2246_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(0)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(0)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*0+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*0)"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(1)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(1)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*1+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*1)"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1010101010101010),
    .INIT_LUTG1(16'b0011000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2249|_al_u2248  (
    .a({open_n12359,_al_u2247_o}),
    .b({_al_u2246_o,\t/a/alu/n145_lutinv }),
    .c({_al_u2161_o,\t/a/alu/n143_lutinv }),
    .d({_al_u2248_o,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 ,\t/a/EX_B [2]}),
    .f({_al_u2249_o,_al_u2248_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2250 (
    .a({\t/a/alu/n5 [28],\t/a/alu/n5 [28]}),
    .b({_al_u2243_o,_al_u2243_o}),
    .c({_al_u2249_o,_al_u2249_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n12394,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .fx({open_n12399,_al_u2250_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1101100011011000),
    .MODE("LOGIC"))
    \_al_u2251|_al_u2257  (
    .a({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [28]}),
    .b({\t/a/EX_A [29],\t/a/EX_B [28]}),
    .c({\t/a/EX_A [28],_al_u2169_o}),
    .d({open_n12404,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .f({\t/a/alu/n19_lutinv ,_al_u2257_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*~C*D+~A*B*~C*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    .INIT_LUTF0(16'b1111010111110101),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0000010100000101),
    .INIT_LUTG1(16'b0000111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2252|_al_u2286  (
    .a({\t/a/alu/n19_lutinv ,\t/a/alu/n21_lutinv }),
    .c({\t/a/alu/n17_lutinv ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/alu/n19_lutinv }),
    .f({_al_u2252_o,_al_u2286_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*A)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(~C*A)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000101000001010),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000101000001010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2253|_al_u2254  (
    .a({open_n12449,\t/a/alu/n104_lutinv }),
    .c({open_n12452,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }),
    .d({_al_u2252_o,open_n12455}),
    .e({\t/a/EX_B [2],open_n12456}),
    .f({\t/a/alu/n104_lutinv ,\t/a/alu/n136_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(A*~(C*B)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000011010101),
    .MODE("LOGIC"))
    \_al_u2256|_al_u2255  (
    .a({_al_u2255_o,\t/a/EX_A [28]}),
    .b({\t/a/alu/n136_lutinv ,\t/a/EX_B [28]}),
    .c({_al_u2161_o,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2256_o,_al_u2255_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*~D*~C+B*~A*~D*~C+~B*~A*D*~C+B*~A*D*~C+~B*~A*~D*C+B*~A*~D*C+~B*~A*D*C+B*~A*D*C"),
    //.LUTF1("~A*~D*~C*~B+~A*~D*C*~B+~A*~D*~C*B+~A*~D*C*B"),
    //.LUTG0("~B*~A*D*~C+B*~A*D*~C+~B*~A*D*C+B*~A*D*C"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*~D*C*B+A*~D*C*B"),
    .INIT_LUTF0(16'b0101010101010101),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b0101010100000000),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2259|_al_u2330  (
    .a({\t/a/alu/n6 [27],_al_u2128_o}),
    .d({_al_u2128_o,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .e({\t/a/EX_operation$0$_lutinv_placeOpt_4 ,\t/a/alu/n6 [23]}),
    .f({_al_u2259_o,_al_u2330_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~D*~C)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~D*~C)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2261|_al_u2379  (
    .c({_al_u2143_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }),
    .d({\t/a/EX_B [2],\t/a/alu/n232_lutinv }),
    .f({\t/a/alu/n232_lutinv ,\t/a/alu/n264_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*B*~D+~A*C*B*~D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTF1("~(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D)"),
    //.LUTG0("~A*~C*B*~D+~A*C*B*~D"),
    //.LUTG1("~(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D)"),
    .INIT_LUTF0(16'b1100110001000100),
    .INIT_LUTF1(16'b0011001110101010),
    .INIT_LUTG0(16'b0000000001000100),
    .INIT_LUTG1(16'b0011001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2262|_al_u2378  (
    .a({_al_u2260_o,_al_u2265_o}),
    .b({\t/a/alu/n232_lutinv ,_al_u2161_o}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }),
    .e({open_n12555,_al_u2260_o}),
    .f({_al_u2262_o,_al_u2378_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~D*~C+A*B*~D*~C+~A*B*D*~C+A*B*D*~C+A*~B*~D*C+A*B*~D*C+A*~B*D*C+A*B*D*C"),
    //.LUTF1("~A*~C*B*~D+~A*C*B*~D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG0("0"),
    //.LUTG1("~A*~C*B*~D+~A*C*B*~D"),
    .INIT_LUTF0(16'b1010110010101100),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2266|_al_u2264  (
    .a({_al_u2264_o,_al_u2150_o}),
    .b({_al_u2161_o,_al_u2157_o}),
    .c({open_n12576,\t/a/EX_B [2]}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 ,open_n12579}),
    .e({_al_u2265_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 }),
    .f({_al_u2266_o,_al_u2264_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2267 (
    .a({\t/a/alu/n5 [27],\t/a/alu/n5 [27]}),
    .b({_al_u2263_o,_al_u2263_o}),
    .c({_al_u2266_o,_al_u2266_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n12612,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .fx({open_n12617,_al_u2267_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    //.LUT1("~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    .INIT_LUT0(16'b1010110010101100),
    .INIT_LUT1(16'b0001000110111011),
    .MODE("LOGIC"))
    \_al_u2269|_al_u2268  (
    .a({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [28]}),
    .b({\t/a/alu/n20_lutinv ,\t/a/EX_A [27]}),
    .c({open_n12620,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n18_lutinv ,open_n12623}),
    .f({_al_u2269_o,\t/a/alu/n20_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUT1("(~D*~C)"),
    .INIT_LUT0(16'b1111101001010000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u2271|_al_u2385  (
    .a({open_n12642,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_1 }),
    .c({_al_u2270_o,_al_u2384_o}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_1 ,_al_u2270_o}),
    .f({\t/a/alu/n135_lutinv ,_al_u2385_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(A*~(C*B)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000011010101),
    .MODE("LOGIC"))
    \_al_u2273|_al_u2272  (
    .a({_al_u2272_o,\t/a/EX_A [27]}),
    .b({\t/a/alu/n135_lutinv ,\t/a/EX_B [27]}),
    .c({_al_u2161_o,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2273_o,_al_u2272_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~C*~A*~D+B*~C*~A*~D+~B*~C*A*~D+B*~C*A*~D+~B*~C*~A*D+B*~C*~A*D+~B*~C*A*D+B*~C*A*D"),
    //.LUTF1("(~C*~(~A*D))"),
    //.LUTG0("~B*~C*A*~D+B*~C*A*~D+~B*~C*A*D+B*~C*A*D"),
    //.LUTG1("(~C*~(~A*D))"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000101000001111),
    .INIT_LUTG0(16'b0000101000001010),
    .INIT_LUTG1(16'b0000101000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2276|_al_u2310  (
    .a({\t/a/EX_operation$0$_lutinv_placeOpt_4 ,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .c({_al_u2128_o,_al_u2128_o}),
    .d({\t/a/alu/n6 [26],open_n12689}),
    .e({open_n12690,\t/a/alu/n6 [24]}),
    .f({_al_u2276_o,_al_u2310_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*D)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTG0("(~A*D)"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0101010100000000),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0101010100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2278|_al_u2391  (
    .a({open_n12711,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_B [2],open_n12714}),
    .d({open_n12717,\t/a/alu/n233_lutinv }),
    .e({_al_u2185_o,open_n12718}),
    .f({\t/a/alu/n233_lutinv ,\t/a/alu/n265_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("~(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0101010111110000),
    .MODE("LOGIC"))
    \_al_u2279|_al_u2390  (
    .a({\t/a/alu/n233_lutinv ,_al_u2282_o}),
    .b({open_n12739,_al_u2277_o}),
    .c({_al_u2277_o,_al_u2161_o}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2279_o,_al_u2390_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~A*~(~0*B))"),
    //.LUTF1("~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG0("(D*~C*~A*~(~1*B))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b1010101010101010),
    .INIT_LUTG0(16'b0000010100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2280|_al_u2284  (
    .a({_al_u2146_o,_al_u2280_o}),
    .b({open_n12760,\t/a/alu/n5 [26]}),
    .c({open_n12761,_al_u2283_o}),
    .d({open_n12764,_al_u2128_o}),
    .e({_al_u2279_o,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .f({_al_u2280_o,_al_u2284_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u2283|_al_u2281  (
    .a({_al_u2281_o,_al_u2198_o}),
    .b({_al_u2282_o,_al_u2191_o}),
    .c({_al_u2161_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .f({_al_u2283_o,_al_u2281_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*C*~A+D*B*C*~A"),
    //.LUTF1("~A*C*~B*D+A*C*~B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*B*C*A+D*B*C*A"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*C*~B*D+A*C*~B*D+~A*C*B*D+A*C*B*D"),
    .INIT_LUTF0(16'b0100000001000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1101000011010000),
    .INIT_LUTG1(16'b1111000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2285|_al_u2291  (
    .a({open_n12805,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .b({open_n12806,\t/a/EX_B [26]}),
    .c({\t/a/EX_A [27],_al_u2169_o}),
    .d({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,open_n12809}),
    .e({\t/a/EX_A [26],\t/a/EX_A [26]}),
    .f({\t/a/alu/n21_lutinv ,_al_u2291_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    //.LUT1("(~A*~B)"),
    .INIT_LUT0(16'b1100101011001010),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"))
    \_al_u2288|_al_u2397  (
    .a({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 ,_al_u2396_o}),
    .b({_al_u2287_o,_al_u2287_o}),
    .c({open_n12830,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }),
    .f({\t/a/alu/n134_lutinv ,_al_u2397_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    //.LUTG0("~B*A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b1111010100000000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b1111101000000000),
    .INIT_LUTG1(16'b0010001000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2290|_al_u2289  (
    .a({\t/a/alu/n134_lutinv ,\t/a/EX_B [26]}),
    .b({\t/a/EX_operation [1],open_n12853}),
    .c({open_n12854,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .d({_al_u2289_o,\t/a/EX_operation [2]}),
    .e({_al_u2161_o,\t/a/EX_A [26]}),
    .f({_al_u2290_o,_al_u2289_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*D)"),
    //.LUT1("(~B*D)"),
    .INIT_LUT0(16'b0101010100000000),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"))
    \_al_u2295|_al_u2402  (
    .a({open_n12877,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_3 }),
    .b({\t/a/EX_B [2],open_n12878}),
    .d({\t/a/alu/n202_lutinv ,\t/a/alu/n234_lutinv }),
    .f({\t/a/alu/n234_lutinv ,\t/a/alu/n266_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*A*D+C*~B*A*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~C*~B*A*D+C*~B*A*D"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b1100110011001100),
    .INIT_LUTG0(16'b0010001000000000),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2296|_al_u2404  (
    .a({\t/a/alu/n234_lutinv ,_al_u2161_o}),
    .b({_al_u2294_o,_al_u2294_o}),
    .d({open_n12905,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_3 }),
    .e({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_3 ,_al_u2299_o}),
    .f({_al_u2296_o,_al_u2404_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~C*~D*~(~0*A))"),
    //.LUTF1("(A*~B)"),
    //.LUTG0("(B*~C*~D*~(~1*A))"),
    //.LUTG1("(A*~B)"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b0010001000100010),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0010001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2297|_al_u2301  (
    .a({_al_u2146_o,\t/a/alu/n5 [25]}),
    .b({_al_u2296_o,_al_u2128_o}),
    .c({open_n12926,_al_u2300_o}),
    .d({open_n12929,_al_u2297_o}),
    .e({open_n12930,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .f({_al_u2297_o,_al_u2301_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(B*~A*~(D*C))"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b0000010001000100),
    .MODE("LOGIC"))
    \_al_u2300|_al_u2298  (
    .a({_al_u2298_o,_al_u2224_o}),
    .b({_al_u2161_o,_al_u2221_o}),
    .c({_al_u2299_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 }),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 ,\t/a/EX_B [2]}),
    .f({_al_u2300_o,_al_u2298_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    //.LUT1("~(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)"),
    .INIT_LUT0(16'b1111101000001010),
    .INIT_LUT1(16'b0100010001110111),
    .MODE("LOGIC"))
    \_al_u2303|_al_u2302  (
    .a({\t/a/alu/n20_lutinv ,\t/a/EX_A [25]}),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n12971}),
    .c({open_n12972,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n22_lutinv ,\t/a/EX_A [26]}),
    .f({_al_u2303_o,\t/a/alu/n22_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2304|_al_u2305  (
    .b({_al_u2229_o,open_n12995}),
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 }),
    .d({_al_u2303_o,_al_u2304_o}),
    .f({_al_u2304_o,\t/a/alu/n133_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(A*~(~C*(B@D)))"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1010100010100010),
    .MODE("LOGIC"))
    \_al_u2306|_al_u1344  (
    .a({\t/a/EX_operation [2],\t/a/ID_rs2$0$_placeOpt_19 }),
    .b({\t/a/EX_B [25],\t/a/ID_rs2$1$_placeOpt_19 }),
    .c({\t/a/EX_operation$0$_lutinv_placeOpt_4 ,\t/a/regfile/regfile$4$ [25]}),
    .d({\t/a/EX_A [25],\t/a/regfile/regfile$5$ [25]}),
    .f({_al_u2306_o,_al_u1344_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~A)"),
    //.LUT1("(~D*~(B*~(C*A)))"),
    .INIT_LUT0(16'b0100010001000100),
    .INIT_LUT1(16'b0000000010110011),
    .MODE("LOGIC"))
    \_al_u2307|_al_u2431  (
    .a({\t/a/alu/n133_lutinv ,\t/a/EX_operation [1]}),
    .b({_al_u2306_o,\t/a/EX_operation [2]}),
    .c({_al_u2161_o,open_n13036}),
    .d({\t/a/EX_operation [1],open_n13039}),
    .f({_al_u2307_o,_al_u2431_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~((~0*~D*B))*~(C)+~A*(~0*~D*B)*~(C)+~(~A)*(~0*~D*B)*C+~A*(~0*~D*B)*C)"),
    //.LUTF1("~A*B*~D*~C+A*B*~D*~C+A*~B*D*~C+A*B*D*~C+~A*B*~D*C+A*B*~D*C+A*~B*D*C+A*B*D*C"),
    //.LUTG0("~(~A*~((~1*~D*B))*~(C)+~A*(~1*~D*B)*~(C)+~(~A)*(~1*~D*B)*C+~A*(~1*~D*B)*C)"),
    //.LUTG1("~A*B*~D*~C+A*B*~D*~C+A*~B*D*~C+A*B*D*~C+~A*B*~D*C+A*B*~D*C+A*~B*D*C+A*B*D*C"),
    .INIT_LUTF0(16'b1111101000111010),
    .INIT_LUTF1(16'b1010101011001100),
    .INIT_LUTG0(16'b1111101011111010),
    .INIT_LUTG1(16'b1010101011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2311|_al_u2312  (
    .a({_al_u2240_o,_al_u2311_o}),
    .b({_al_u2238_o,_al_u2184_o}),
    .c({open_n13058,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_B [2],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({open_n13061,\t/a/EX_B [2]}),
    .f({_al_u2311_o,_al_u2312_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b1111101000001010),
    .MODE("LOGIC"))
    \_al_u2315|_al_u2415  (
    .a({_al_u2245_o,_al_u2315_o}),
    .b({open_n13082,_al_u2311_o}),
    .c({\t/a/EX_B [2],_al_u2161_o}),
    .d({_al_u2237_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_1 }),
    .f({_al_u2315_o,_al_u2415_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("0"),
    //.LUTG1("~A*~B*C*~D+~A*~B*C*D"),
    .INIT_LUTF0(16'b1100110010101010),
    .INIT_LUTF1(16'b0101000001010000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0001000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2316|_al_u2314  (
    .a({_al_u2314_o,_al_u2247_o}),
    .b({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 ,_al_u2244_o}),
    .c({_al_u2161_o,open_n13103}),
    .d({open_n13106,\t/a/EX_B [2]}),
    .e({_al_u2315_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 }),
    .f({_al_u2316_o,_al_u2314_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2317 (
    .a({\t/a/alu/n5 [24],\t/a/alu/n5 [24]}),
    .b({_al_u2313_o,_al_u2313_o}),
    .c({_al_u2316_o,_al_u2316_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n13139,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .fx({open_n13144,_al_u2317_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1101110110001000),
    .MODE("LOGIC"))
    \_al_u2318|_al_u2324  (
    .a({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [24]}),
    .b({\t/a/EX_A [25],\t/a/EX_B [24]}),
    .c({open_n13147,_al_u2169_o}),
    .d({\t/a/EX_A [24],\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .f({\t/a/alu/n23_lutinv ,_al_u2324_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    //.LUTG1("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0101111101011111),
    .INIT_LUTF1(16'b0101111101011111),
    .INIT_LUTG0(16'b0101000001010000),
    .INIT_LUTG1(16'b0101000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2319|_al_u2345  (
    .a({\t/a/alu/n21_lutinv ,\t/a/alu/n23_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/alu/n23_lutinv ,\t/a/alu/n25_lutinv }),
    .f({_al_u2319_o,_al_u2345_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    //.LUTF1("~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG0("~D*~C*~B*~A+D*~C*~B*~A+~D*C*~B*~A+D*C*~B*~A+~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+D*C*~B*A+~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    //.LUTG1("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    .INIT_LUTF0(16'b1000100010001000),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b1011101110111011),
    .INIT_LUTG1(16'b1111111101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2320|_al_u2372  (
    .a({\t/a/EX_B [2],_al_u2319_o}),
    .b({open_n13194,\t/a/EX_B [2]}),
    .d({_al_u2252_o,open_n13199}),
    .e({_al_u2319_o,_al_u2371_o}),
    .f({_al_u2320_o,_al_u2372_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    //.LUTF1("(~A*~D)"),
    //.LUTG0("(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    //.LUTG1("(~A*~D)"),
    .INIT_LUTF0(16'b1110111000100010),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b1110111000100010),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2321|_al_u2422  (
    .a({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,_al_u2421_o}),
    .b({open_n13220,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2320_o,_al_u2320_o}),
    .f({\t/a/alu/n132_lutinv ,_al_u2422_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*~A*C+~B*D*~A*C+~B*~D*A*C+B*~D*A*C+~B*D*A*C+B*D*A*C"),
    //.LUTF1("~A*~B*~D*~C+~A*~B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    //.LUTG0("B*~D*~A*C+B*D*~A*C+~B*~D*A*C+B*~D*A*C+~B*D*A*C+B*D*A*C"),
    //.LUTG1("~A*~B*~D*~C+~A*~B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*~B*D*C+A*~B*D*C"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b1110000011100000),
    .INIT_LUTG1(16'b0011000100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2323|_al_u2322  (
    .a({_al_u2322_o,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .b({\t/a/EX_operation [1],\t/a/EX_A [24]}),
    .c({\t/a/alu/n132_lutinv ,\t/a/EX_operation [2]}),
    .e({_al_u2161_o,\t/a/EX_B [24]}),
    .f({_al_u2323_o,_al_u2322_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D)"),
    //.LUT1("(~D*~C)"),
    .INIT_LUT0(16'b1111000010101010),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u2326|_al_u2145  (
    .a({open_n13271,_al_u2137_o}),
    .c({_al_u2144_o,_al_u2144_o}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({\t/a/alu/n260_lutinv ,_al_u2145_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("0"),
    //.LUTG0("0"),
    //.LUTG1("~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2327|_al_u2540  (
    .a({_al_u2146_o,_al_u2128_o}),
    .e({\t/a/alu/n260_lutinv ,_al_u2539_o}),
    .f({_al_u2327_o,_al_u2540_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2329 (
    .a({\t/a/alu/n5 [23],\t/a/alu/n5 [23]}),
    .b({_al_u2327_o,_al_u2327_o}),
    .c({_al_u2328_o,_al_u2328_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n13334,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .fx({open_n13339,_al_u2329_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~D*~C+A*B*~D*~C+A*~B*D*~C+A*B*D*~C+A*~B*~D*C+A*B*~D*C+A*~B*D*C+A*B*D*C"),
    //.LUTF1("~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)"),
    //.LUTG0("~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG1("~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0011001101010101),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0011001101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2332|_al_u2331  (
    .a({\t/a/alu/n24_lutinv ,\t/a/EX_A [23]}),
    .b({\t/a/alu/n22_lutinv ,open_n13342}),
    .c({open_n13343,\t/a/EX_A [24]}),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n13346}),
    .e({open_n13347,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2332_o,\t/a/alu/n24_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~C*~D*~B+A*C*~D*~B+A*~C*D*~B+A*C*D*~B+A*~C*~D*B+A*C*~D*B+A*~C*D*B+A*C*D*B"),
    //.LUTF1("~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    //.LUTG0("~A*~C*~D*~B+A*~C*~D*~B+~A*~C*D*~B+A*~C*D*~B+~A*~C*~D*B+A*~C*~D*B+~A*C*~D*B+A*C*~D*B+~A*~C*D*B+A*~C*D*B+~A*C*D*B+A*C*D*B"),
    //.LUTG1("~D*~C*~B*~A+D*~C*~B*~A+~D*C*~B*~A+D*C*~B*~A+~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+D*C*~B*A+~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1100111111001111),
    .INIT_LUTG1(16'b1011101110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2333|_al_u2334  (
    .a({_al_u2269_o,_al_u2333_o}),
    .b({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .c({open_n13368,\t/a/alu/n56_lutinv }),
    .e({_al_u2332_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2333_o,_al_u2334_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(A*~(C*~B)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000001110101),
    .MODE("LOGIC"))
    \_al_u2336|_al_u2335  (
    .a({_al_u2335_o,\t/a/EX_A [23]}),
    .b({_al_u2334_o,\t/a/EX_B [23]}),
    .c({_al_u2161_o,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2336_o,_al_u2335_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    //.LUTF1("(~C*~A)"),
    //.LUTG0("(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    //.LUTG1("(~C*~A)"),
    .INIT_LUTF0(16'b1010111110100000),
    .INIT_LUTF1(16'b0000010100000101),
    .INIT_LUTG0(16'b1010111110100000),
    .INIT_LUTG1(16'b0000010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2339|_al_u2187  (
    .a({_al_u2186_o,_al_u2186_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }),
    .d({open_n13417,_al_u2179_o}),
    .f({\t/a/alu/n261_lutinv ,_al_u2187_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~C*~D*~(~0*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*~C*~D*~(~1*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000000100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2340|_al_u2342  (
    .a({open_n13440,\t/a/alu/n5 [22]}),
    .b({open_n13441,_al_u2128_o}),
    .c({_al_u2146_o,_al_u2341_o}),
    .d({\t/a/alu/n261_lutinv ,_al_u2340_o}),
    .e({open_n13444,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .f({_al_u2340_o,_al_u2342_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1111000010101010),
    .MODE("LOGIC"))
    \_al_u2344|_al_u2350  (
    .a({\t/a/EX_A [22],\t/a/EX_A [22]}),
    .b({open_n13465,\t/a/EX_B [22]}),
    .c({\t/a/EX_A [23],_al_u2169_o}),
    .d({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .f({\t/a/alu/n25_lutinv ,_al_u2350_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    //.LUT1("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    .INIT_LUT0(16'b1110111001000100),
    .INIT_LUT1(16'b1110111001000100),
    .MODE("LOGIC"))
    \_al_u2346|_al_u2396  (
    .a({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .b({_al_u2345_o,_al_u2395_o}),
    .d({_al_u2286_o,_al_u2345_o}),
    .f({_al_u2346_o,_al_u2396_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(A*~(C*~B)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000001110101),
    .MODE("LOGIC"))
    \_al_u2349|_al_u2348  (
    .a({_al_u2348_o,\t/a/EX_A [22]}),
    .b({_al_u2347_o,\t/a/EX_B [22]}),
    .c({_al_u2161_o,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2349_o,_al_u2348_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A)"),
    //.LUT1("(~A*~B)"),
    .INIT_LUT0(16'b1101110110001000),
    .INIT_LUT1(16'b0001000100010001),
    .MODE("LOGIC"))
    \_al_u2352|_al_u2219  (
    .a({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 }),
    .b({_al_u2218_o,_al_u2218_o}),
    .d({open_n13532,_al_u2215_o}),
    .f({\t/a/alu/n262_lutinv ,_al_u2219_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~A*~(~0*B))"),
    //.LUTF1("(B*D)"),
    //.LUTG0("(D*~C*~A*~(~1*B))"),
    //.LUTG1("(B*D)"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b1100110000000000),
    .INIT_LUTG0(16'b0000010100000000),
    .INIT_LUTG1(16'b1100110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2353|_al_u2355  (
    .a({open_n13551,_al_u2353_o}),
    .b({_al_u2146_o,\t/a/alu/n5 [21]}),
    .c({open_n13552,_al_u2354_o}),
    .d({\t/a/alu/n262_lutinv ,_al_u2128_o}),
    .e({open_n13555,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .f({_al_u2353_o,_al_u2355_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)"),
    //.LUTG0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0011001101010101),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b0011001101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2358|_al_u2357  (
    .a({\t/a/alu/n26_lutinv ,\t/a/EX_A [21]}),
    .b({\t/a/alu/n24_lutinv ,open_n13576}),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [22]}),
    .e({open_n13581,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2358_o,\t/a/alu/n26_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*D*A+C*~B*D*A+~C*B*D*A+C*B*D*A"),
    //.LUTF1("A*~B*D*~C+A*B*D*~C+A*~B*D*C+A*B*D*C"),
    //.LUTG0("~C*~B*~D*~A+C*~B*~D*~A+~C*B*~D*~A+C*B*~D*~A+~C*~B*~D*A+C*~B*~D*A+~C*B*~D*A+C*B*~D*A+~C*~B*D*A+C*~B*D*A+~C*B*D*A+C*B*D*A"),
    //.LUTG1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+A*~B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+A*~B*D*C+A*B*D*C"),
    .INIT_LUTF0(16'b1010101000000000),
    .INIT_LUTF1(16'b1010101000000000),
    .INIT_LUTG0(16'b1010101011111111),
    .INIT_LUTG1(16'b1010101011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2359|_al_u2409  (
    .a({_al_u2303_o,_al_u2358_o}),
    .d({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .e({_al_u2358_o,_al_u2408_o}),
    .f({_al_u2359_o,_al_u2409_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*~A*C+~B*D*~A*C+~B*~D*A*C+B*~D*A*C+~B*D*A*C+B*D*A*C"),
    //.LUTF1("~B*~A*~C*~D+~B*A*~C*~D+~B*~A*C*~D+~B*A*C*~D+~B*~A*C*D+~B*A*C*D"),
    //.LUTG0("B*~D*~A*C+B*D*~A*C+~B*~D*A*C+B*~D*A*C+~B*D*A*C+B*D*A*C"),
    //.LUTG1("~B*~A*~C*~D+~B*A*~C*~D+~B*~A*C*~D+~B*A*C*~D"),
    .INIT_LUTF0(16'b1011000010110000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b1110000011100000),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2362|_al_u2361  (
    .a({open_n13628,\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .b({\t/a/EX_operation [1],\t/a/EX_A [21]}),
    .c({_al_u2161_o,\t/a/EX_operation [2]}),
    .d({_al_u2361_o,open_n13631}),
    .e({_al_u2360_o,\t/a/EX_B [21]}),
    .f({_al_u2362_o,_al_u2361_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~D)"),
    //.LUT1("(D*A)"),
    .INIT_LUT0(16'b0000000000110011),
    .INIT_LUT1(16'b1010101000000000),
    .MODE("LOGIC"))
    \_al_u2366|_al_u2365  (
    .a({\t/a/alu/n263_lutinv ,open_n13652}),
    .b({open_n13653,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2146_o,_al_u2241_o}),
    .f({_al_u2366_o,\t/a/alu/n263_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2368 (
    .a({\t/a/alu/n5 [20],\t/a/alu/n5 [20]}),
    .b({_al_u2366_o,_al_u2366_o}),
    .c({_al_u2367_o,_al_u2367_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n13688,\t/a/EX_operation$0$_lutinv_placeOpt_2 }),
    .fx({open_n13693,_al_u2368_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1110111000100010),
    .MODE("LOGIC"))
    \_al_u2370|_al_u2376  (
    .a({\t/a/EX_A [20],\t/a/EX_A [20]}),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [20]}),
    .c({open_n13696,_al_u2169_o}),
    .d({\t/a/EX_A [21],\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .f({\t/a/alu/n27_lutinv ,_al_u2376_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0100010001110111),
    .MODE("LOGIC"))
    \_al_u2371|_al_u2395  (
    .a({\t/a/alu/n25_lutinv ,open_n13717}),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/alu/n29_lutinv }),
    .c({open_n13718,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n27_lutinv ,\t/a/alu/n27_lutinv }),
    .f({_al_u2371_o,_al_u2395_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~D*~B+A*~C*~D*~B+~A*~C*D*~B+A*~C*D*~B"),
    //.LUTF1("~(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)"),
    //.LUTG0("~A*~C*~D*~B+A*~C*~D*~B+~A*C*~D*~B+~A*~C*D*~B+A*~C*D*~B+~A*C*D*~B"),
    //.LUTG1("~(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D)"),
    .INIT_LUTF0(16'b0000001100000011),
    .INIT_LUTF1(16'b0101010111110000),
    .INIT_LUTG0(16'b0001001100010011),
    .INIT_LUTG1(16'b0101010111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2373|_al_u2375  (
    .a({\t/a/alu/n104_lutinv ,_al_u2373_o}),
    .b({open_n13739,\t/a/EX_operation [1]}),
    .c({_al_u2372_o,_al_u2374_o}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 ,open_n13742}),
    .e({open_n13743,_al_u2161_o}),
    .f({_al_u2373_o,_al_u2375_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*~C*~A+D*~B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+D*~B*C*A"),
    //.LUTF1("0"),
    //.LUTG0("~D*~B*~C*~A+~D*~B*~C*A"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b1111101011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2374|_al_u743  (
    .a({\t/a/EX_A [20],open_n13764}),
    .b({open_n13765,\t/a/ID_rs1$1$_placeOpt_15 }),
    .c({\t/a/EX_operation$0$_lutinv_placeOpt_4 ,\t/a/regfile/regfile$4$ [20]}),
    .d({\t/a/EX_B [20],\t/a/ID_rs1$0$_placeOpt_15 }),
    .e({\t/a/EX_operation [2],\t/a/regfile/regfile$5$ [20]}),
    .f({_al_u2374_o,_al_u743_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(A*~((~C*B))*~(0)+A*(~C*B)*~(0)+~(A)*(~C*B)*0+A*(~C*B)*0))"),
    //.LUTF1("(~B*~(A*~((D*C))*~(0)+A*(D*C)*~(0)+~(A)*(D*C)*0+A*(D*C)*0))"),
    //.LUTG0("(~D*(A*~((~C*B))*~(1)+A*(~C*B)*~(1)+~(A)*(~C*B)*1+A*(~C*B)*1))"),
    //.LUTG1("(~B*~(A*~((D*C))*~(1)+A*(D*C)*~(1)+~(A)*(D*C)*1+A*(D*C)*1))"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2380|_al_u2549  (
    .a({\t/a/alu/n5 [19],\t/a/alu/n5 [3]}),
    .b({_al_u2378_o,\t/a/alu/n264_lutinv }),
    .c({\t/a/alu/n264_lutinv ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation [1]}),
    .e({\t/a/EX_operation$0$_lutinv_placeOpt_5 ,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .f({_al_u2380_o,\t/a/alu/mux0_b3/B1_0 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~A*D))"),
    //.LUT1("(~B*~(~C*A))"),
    .INIT_LUT0(16'b0010001000110011),
    .INIT_LUT1(16'b0011000100110001),
    .MODE("LOGIC"))
    \_al_u2381|_al_u2293  (
    .a({\t/a/alu/n6 [19],\t/a/EX_operation$0$_lutinv_placeOpt_4 }),
    .b({\t/a/EX_operation [2],_al_u2128_o}),
    .c({_al_u2128_o,open_n13810}),
    .d({open_n13813,\t/a/alu/n6 [25]}),
    .f({_al_u2381_o,_al_u2293_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    //.LUT1("~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    .INIT_LUT0(16'b1110010011100100),
    .INIT_LUT1(16'b0101000001011111),
    .MODE("LOGIC"))
    \_al_u2383|_al_u2382  (
    .a({\t/a/alu/n26_lutinv ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .b({open_n13832,\t/a/EX_A [19]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [20]}),
    .d({\t/a/alu/n28_lutinv ,open_n13835}),
    .f({_al_u2383_o,\t/a/alu/n28_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*~A*D+C*~B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("~A*~B*~D*~C+~A*~B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    //.LUTG0("~C*B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG1("~A*~B*~D*~C+A*~B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    .INIT_LUTF0(16'b1011101100000000),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b1110111000000000),
    .INIT_LUTG1(16'b0001001100010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2387|_al_u2386  (
    .a({_al_u2386_o,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .b({\t/a/EX_operation [1],\t/a/EX_B [19]}),
    .c({_al_u2385_o,open_n13854}),
    .d({open_n13857,\t/a/EX_operation [2]}),
    .e({_al_u2161_o,\t/a/EX_A [19]}),
    .f({_al_u2387_o,_al_u2386_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(A*~((~C*B))*~(0)+A*(~C*B)*~(0)+~(A)*(~C*B)*0+A*(~C*B)*0))"),
    //.LUTF1("(~B*~(A*~((D*C))*~(0)+A*(D*C)*~(0)+~(A)*(D*C)*0+A*(D*C)*0))"),
    //.LUTG0("(~D*(A*~((~C*B))*~(1)+A*(~C*B)*~(1)+~(A)*(~C*B)*1+A*(~C*B)*1))"),
    //.LUTG1("(~B*~(A*~((D*C))*~(1)+A*(D*C)*~(1)+~(A)*(D*C)*1+A*(D*C)*1))"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2392|_al_u2558  (
    .a({\t/a/alu/n5 [18],\t/a/alu/n5 [2]}),
    .b({_al_u2390_o,\t/a/alu/n265_lutinv }),
    .c({\t/a/alu/n265_lutinv ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation [1]}),
    .e({\t/a/EX_operation$0$_lutinv_placeOpt_1 ,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .f({_al_u2392_o,\t/a/alu/mux0_b2/B1_0 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~B*~(~C*~A)))"),
    //.LUT1("(~C*~(~A*D))"),
    .INIT_LUT0(16'b1100110100000000),
    .INIT_LUT1(16'b0000101000001111),
    .MODE("LOGIC"))
    \_al_u2393|_al_u2728  (
    .a({_al_u2128_o,\t/a/alu/mux0_b6/B1_0 }),
    .b({open_n13900,_al_u2526_o}),
    .c({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .d({\t/a/alu/n6 [18],_al_u2128_o}),
    .f({_al_u2393_o,_al_u2728_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1100101011001010),
    .MODE("LOGIC"))
    \_al_u2394|_al_u2400  (
    .a({\t/a/EX_A [18],\t/a/EX_A [18]}),
    .b({\t/a/EX_A [19],\t/a/EX_B [18]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({open_n13923,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .f({\t/a/alu/n29_lutinv ,_al_u2400_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(A*~(C*~B)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000001110101),
    .MODE("LOGIC"))
    \_al_u2399|_al_u2398  (
    .a({_al_u2398_o,\t/a/EX_A [18]}),
    .b({_al_u2397_o,\t/a/EX_B [18]}),
    .c({_al_u2161_o,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2399_o,_al_u2398_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(A*~((~C*B))*~(0)+A*(~C*B)*~(0)+~(A)*(~C*B)*0+A*(~C*B)*0))"),
    //.LUTF1("(A*B)"),
    //.LUTG0("(~D*(A*~((~C*B))*~(1)+A*(~C*B)*~(1)+~(A)*(~C*B)*1+A*(~C*B)*1))"),
    //.LUTG1("(A*B)"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2403|_al_u2579  (
    .a({_al_u2146_o,\t/a/alu/n5 [1]}),
    .b({\t/a/alu/n266_lutinv ,\t/a/alu/n266_lutinv }),
    .c({open_n13962,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({open_n13965,\t/a/EX_operation [1]}),
    .e({open_n13966,\t/a/EX_operation [0]}),
    .f({_al_u2403_o,\t/a/alu/mux0_b1/B1_0 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2405 (
    .a({\t/a/alu/n5 [17],\t/a/alu/n5 [17]}),
    .b({_al_u2403_o,_al_u2403_o}),
    .c({_al_u2404_o,_al_u2404_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n13999,\t/a/EX_operation [0]}),
    .fx({open_n14004,_al_u2405_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~D*C*~B+A*D*C*~B"),
    //.LUTF1("A*~B*~D*~C+A*B*~D*~C+A*~B*~D*C+A*B*~D*C"),
    //.LUTG0("~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+A*~D*C*B+A*D*C*B"),
    //.LUTG1("A*~B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+A*~B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    .INIT_LUTF0(16'b0010000000100000),
    .INIT_LUTF1(16'b0000000010101010),
    .INIT_LUTG0(16'b1011000010110000),
    .INIT_LUTG1(16'b1111111110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2407|_al_u2413  (
    .a({\t/a/EX_A [17],\t/a/EX_A [17]}),
    .b({open_n14007,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .c({open_n14008,_al_u2169_o}),
    .d({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,open_n14011}),
    .e({\t/a/EX_A [18],\t/a/EX_B [17]}),
    .f({\t/a/alu/n30_lutinv ,_al_u2413_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(B*~(C*~A)))"),
    //.LUT1("(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)"),
    .INIT_LUT0(16'b0000000001110011),
    .INIT_LUT1(16'b1010101011110000),
    .MODE("LOGIC"))
    \_al_u2410|_al_u2412  (
    .a({_al_u2304_o,_al_u2410_o}),
    .b({open_n14032,_al_u2411_o}),
    .c({_al_u2409_o,_al_u2161_o}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 ,\t/a/EX_operation [1]}),
    .f({_al_u2410_o,_al_u2412_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(B*~(~D*(A@C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b1100110010000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2411|t/a/id_ex/reg4_b2  (
    .a({\t/a/EX_B [17],\t/a/aluin/sel1_b17/B9 }),
    .b({\t/a/EX_operation [2],_al_u2007_o}),
    .c({\t/a/EX_A [17],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [0],\t/a/EX_rs1 [2]}),
    .mi({open_n14064,\t/a/ID_rs1$2$_placeOpt_9 }),
    .sr(rst_pad),
    .f({_al_u2411_o,\t/a/EX_B [17]}),
    .q({open_n14068,\t/a/EX_rs1 [2]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*B*A)"),
    //.LUTF1("(D*~(~A*~B*~(~0*C)))"),
    //.LUTG0("(~1*~D*~C*B*A)"),
    //.LUTG1("(D*~(~A*~B*~(~1*C)))"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b1111111000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1110111000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2417|_al_u2416  (
    .a({_al_u2416_o,_al_u2184_o}),
    .b({_al_u2415_o,_al_u2146_o}),
    .c({\t/a/alu/n5 [16],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2128_o,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/EX_operation$0$_lutinv_placeOpt_1 ,\t/a/EX_B [2]}),
    .f({_al_u2417_o,_al_u2416_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*~(D*~A)))"),
    //.LUT1("(~B*~(~C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110110011111100),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2418|t/a/ex_mem/reg4_b16  (
    .a({open_n14091,_al_u2417_o}),
    .b({\t/a/EX_operation [2],_al_u2425_o}),
    .c({_al_u2128_o,_al_u2424_o}),
    .clk(clock_pad),
    .d({\t/a/alu/n6 [16],_al_u2418_o}),
    .sr(rst_pad),
    .f({_al_u2418_o,\t/a/aludat [16]}),
    .q({open_n14108,\t/a/MEM_aludat [16]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0001000111011101),
    .MODE("LOGIC"))
    \_al_u2420|_al_u2419  (
    .a({\t/a/alu/n31_lutinv ,open_n14109}),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [16]}),
    .c({open_n14110,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n29_lutinv ,\t/a/EX_A [17]}),
    .f({_al_u2420_o,\t/a/alu/n31_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111111100001111),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2421|_al_u2463  (
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2420_o,_al_u2420_o}),
    .e({_al_u2371_o,_al_u2462_o}),
    .f({_al_u2421_o,_al_u2463_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(A*~(C*~B)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000001110101),
    .MODE("LOGIC"))
    \_al_u2424|_al_u2423  (
    .a({_al_u2423_o,\t/a/EX_A [16]}),
    .b({_al_u2422_o,\t/a/EX_B [16]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2424_o,_al_u2423_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(A*~((~C*~B))*~(0)+A*(~C*~B)*~(0)+~(A)*(~C*~B)*0+A*(~C*~B)*0))"),
    //.LUT1("(~D*~(A*~((~C*~B))*~(1)+A*(~C*~B)*~(1)+~(A)*(~C*~B)*1+A*(~C*~B)*1))"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2427 (
    .a({\t/a/alu/n5 [15],\t/a/alu/n5 [15]}),
    .b({_al_u2145_o,_al_u2145_o}),
    .c({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n14189,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .fx({open_n14194,_al_u2427_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~C*D*A+B*~C*D*A+~B*C*D*A+B*C*D*A"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A"),
    //.LUTG0("~B*~C*~D*~A+B*~C*~D*~A+~B*C*~D*~A+B*C*~D*~A+~B*~C*~D*A+B*~C*~D*A+~B*C*~D*A+B*C*~D*A+~B*~C*D*A+B*~C*D*A+~B*C*D*A+B*C*D*A"),
    //.LUTG1("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    .INIT_LUTF0(16'b1010101000000000),
    .INIT_LUTF1(16'b0101111101011111),
    .INIT_LUTG0(16'b1010101011111111),
    .INIT_LUTG1(16'b0101000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2429|_al_u2428  (
    .a({\t/a/alu/n30_lutinv ,\t/a/EX_A [16]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n14199}),
    .d({open_n14202,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/alu/n32_lutinv ,\t/a/EX_A [15]}),
    .f({_al_u2429_o,\t/a/alu/n32_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    //.LUT1("(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    .INIT_LUT0(16'b1010111110100000),
    .INIT_LUT1(16'b1010111110100000),
    .MODE("LOGIC"))
    \_al_u2430|_al_u2473  (
    .a({_al_u2383_o,_al_u2429_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2429_o,_al_u2472_o}),
    .f({_al_u2430_o,_al_u2473_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(A*~(~D*(B@C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b1010101010000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2432|t/a/id_ex/reg4_b0  (
    .a({_al_u2431_o,\t/a/aluin/sel1_b15/B9 }),
    .b({\t/a/EX_B [15],_al_u2007_o}),
    .c({\t/a/EX_A [15],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [0],\t/a/EX_rs1 [0]}),
    .mi({open_n14256,\t/a/ID_rs1$0$_placeOpt_20 }),
    .sr(rst_pad),
    .f({_al_u2432_o,\t/a/EX_B [15]}),
    .q({open_n14260,\t/a/EX_rs1 [0]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~D*C*A))"),
    //.LUTF1("(D*~(C*~(A*~(B)*~(0)+A*B*~(0)+~(A)*B*0+A*B*0)))"),
    //.LUTG0("(B*~(~1*~D*C*A))"),
    //.LUTG1("(D*~(C*~(A*~(B)*~(1)+A*B*~(1)+~(A)*B*1+A*B*1)))"),
    .INIT_LUTF0(16'b1100110001001100),
    .INIT_LUTF1(16'b1010111100000000),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2434|_al_u2433  (
    .a({_al_u2430_o,\t/a/alu/n56_lutinv }),
    .b({_al_u2333_o,_al_u2432_o}),
    .c({_al_u2161_o,_al_u2146_o}),
    .d({_al_u2433_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .f({_al_u2434_o,_al_u2433_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~A))"),
    //.LUT1("(~C*~(B*~A))"),
    .INIT_LUT0(16'b0010001000110011),
    .INIT_LUT1(16'b0000101100001011),
    .MODE("LOGIC"))
    \_al_u2435|_al_u2555  (
    .a({\t/a/alu/n6 [15],\t/a/alu/n6 [3]}),
    .b({_al_u2126_o,_al_u2554_o}),
    .c({_al_u2434_o,open_n14283}),
    .d({open_n14286,_al_u2126_o}),
    .f({_al_u2435_o,_al_u2555_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~(~D*A))"),
    //.LUT1("(C*~D*~(~B*A))"),
    .INIT_LUT0(16'b0011000000010000),
    .INIT_LUT1(16'b0000000011010000),
    .MODE("LOGIC"))
    \_al_u2438|_al_u2478  (
    .a({\t/a/alu/n5 [14],\t/a/alu/n5 [10]}),
    .b({\t/a/EX_operation$0$_lutinv_placeOpt_2 ,\t/a/EX_operation [2]}),
    .c({_al_u2128_o,_al_u2128_o}),
    .d({\t/a/EX_operation [2],\t/a/EX_operation$0$_lutinv_placeOpt_2 }),
    .f({_al_u2438_o,_al_u2478_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+D*~B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+D*~B*C*A+D*B*C*A"),
    //.LUTG0("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0001000011110000),
    .INIT_LUTF1(16'b1111111100001111),
    .INIT_LUTG0(16'b0111000011110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2440|_al_u2439  (
    .a({open_n14325,\t/a/EX_A [14]}),
    .b({open_n14326,\t/a/EX_B [14]}),
    .c({_al_u2126_o,\t/a/EX_operation [1]}),
    .d({\t/a/alu/n6 [14],\t/a/EX_operation [2]}),
    .e({_al_u2439_o,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .f({_al_u2440_o,_al_u2439_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*D*~B*~A+C*D*~B*~A+~C*D*~B*A+C*D*~B*A"),
    //.LUTF1("~D*~B*~A*~C+~D*B*~A*~C+~D*~B*A*~C+D*~B*A*~C+~D*B*A*~C+D*B*A*~C+~D*~B*~A*C+~D*B*~A*C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTG0("~C*D*~B*~A+C*D*~B*~A+~C*~D*B*~A+C*~D*B*~A+~C*D*B*~A+C*D*B*~A+~C*D*~B*A+C*D*~B*A+~C*~D*B*A+C*~D*B*A+~C*D*B*A+C*D*B*A"),
    //.LUTG1("~D*~B*~A*~C+~D*B*~A*~C+~D*~B*~A*C+~D*B*~A*C"),
    .INIT_LUTF0(16'b0011001100000000),
    .INIT_LUTF1(16'b1010101011111111),
    .INIT_LUTG0(16'b1111111111001100),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2442|_al_u2441  (
    .a({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n14349}),
    .b({open_n14350,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n33_lutinv ,\t/a/EX_A [14]}),
    .e({\t/a/alu/n31_lutinv ,\t/a/EX_A [15]}),
    .f({_al_u2442_o,\t/a/alu/n33_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    //.LUT1("(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B)"),
    .INIT_LUT0(16'b1110111001000100),
    .INIT_LUT1(16'b1011101110001000),
    .MODE("LOGIC"))
    \_al_u2443|_al_u2483  (
    .a({_al_u2395_o,\t/a/EX_B [2]}),
    .b({\t/a/EX_B [2],_al_u2482_o}),
    .d({_al_u2442_o,_al_u2442_o}),
    .f({_al_u2443_o,_al_u2483_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*~D+C*~B*A*~D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("0"),
    //.LUTG0("~C*~B*A*~D+C*~B*A*~D"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000100010),
    .INIT_LUTG1(16'b0000000001011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2446|_al_u2444  (
    .a({\t/a/alu/n138_lutinv ,_al_u2161_o}),
    .b({open_n14397,_al_u2443_o}),
    .c({_al_u2146_o,open_n14398}),
    .d({_al_u2444_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }),
    .e({_al_u2445_o,_al_u2346_o}),
    .f({_al_u2446_o,_al_u2444_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~(~D*A))"),
    //.LUT1("(C*~B*~(~D*A))"),
    .INIT_LUT0(16'b0011000000010000),
    .INIT_LUT1(16'b0011000000010000),
    .MODE("LOGIC"))
    \_al_u2448|_al_u2508  (
    .a({\t/a/alu/n5 [13],\t/a/alu/n5 [7]}),
    .b({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .c({_al_u2128_o,_al_u2128_o}),
    .d({\t/a/EX_operation$0$_lutinv_placeOpt_1 ,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .f({_al_u2448_o,_al_u2508_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUTF1("(~A*~(B*~D))"),
    //.LUTG0("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    //.LUTG1("(~A*~(B*~D))"),
    .INIT_LUTF0(16'b0001000011110000),
    .INIT_LUTF1(16'b0101010100010001),
    .INIT_LUTG0(16'b0111000011110000),
    .INIT_LUTG1(16'b0101010100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2450|_al_u2449  (
    .a({_al_u2449_o,\t/a/EX_A [13]}),
    .b({_al_u2126_o,\t/a/EX_B [13]}),
    .c({open_n14441,\t/a/EX_operation [1]}),
    .d({\t/a/alu/n6 [13],\t/a/EX_operation [2]}),
    .e({open_n14444,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .f({_al_u2450_o,_al_u2449_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    //.LUT1("~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    .INIT_LUT0(16'b1010101011001100),
    .INIT_LUT1(16'b0101000001011111),
    .MODE("LOGIC"))
    \_al_u2452|_al_u2451  (
    .a({\t/a/alu/n32_lutinv ,\t/a/EX_A [14]}),
    .b({open_n14465,\t/a/EX_A [13]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n14466}),
    .d({\t/a/alu/n34_lutinv ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2452_o,\t/a/alu/n34_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("~C*A*B*~D+C*A*B*~D+~C*A*B*D+C*A*B*D"),
    //.LUTG0("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG1("~C*~A*~B*~D+C*~A*~B*~D+~C*A*~B*~D+C*A*~B*~D+~C*A*B*~D+C*A*B*~D+~C*~A*~B*D+C*~A*~B*D+~C*A*~B*D+C*A*~B*D+~C*A*B*D+C*A*B*D"),
    .INIT_LUTF0(16'b1010101000000000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1111111101010101),
    .INIT_LUTG1(16'b1011101110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2453|_al_u2493  (
    .a({_al_u2408_o,\t/a/EX_B [2]}),
    .b({\t/a/EX_B [2],open_n14487}),
    .d({open_n14492,_al_u2452_o}),
    .e({_al_u2452_o,_al_u2492_o}),
    .f({_al_u2453_o,_al_u2493_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    .INIT_LUTF0(16'b0101000011110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0101000000000000),
    .INIT_LUTG1(16'b0001000101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2456|_al_u2454  (
    .a({_al_u2454_o,_al_u2359_o}),
    .b({\t/a/alu/n137_lutinv ,open_n14513}),
    .c({open_n14514,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 }),
    .e({_al_u2455_o,_al_u2453_o}),
    .f({_al_u2456_o,_al_u2454_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~C*D*~A+B*~C*D*~A+~B*~C*D*A+B*~C*D*A"),
    //.LUTF1("~A*~C*D*~B+~A*~C*D*B"),
    //.LUTG0("~B*~C*D*A+B*~C*D*A"),
    //.LUTG1("~A*~C*D*~B+A*~C*D*~B+~A*~C*D*B+A*~C*D*B"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000010100000000),
    .INIT_LUTG0(16'b0000101000000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2458|_al_u2498  (
    .a({\t/a/alu/n5 [12],\t/a/EX_operation$0$_lutinv_placeOpt_2 }),
    .c({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .d({_al_u2128_o,_al_u2128_o}),
    .e({\t/a/EX_operation$0$_lutinv_placeOpt_2 ,\t/a/alu/n5 [8]}),
    .f({_al_u2458_o,_al_u2498_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUT1("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    .INIT_LUT0(16'b0001000011110000),
    .INIT_LUT1(16'b0111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2459 (
    .a({\t/a/EX_A [12],\t/a/EX_A [12]}),
    .b({\t/a/EX_B [12],\t/a/EX_B [12]}),
    .c({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n14573,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .fx({open_n14578,_al_u2459_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(C*~B))"),
    //.LUT1("(~A*~(C*~D))"),
    .INIT_LUT0(16'b0100010101000101),
    .INIT_LUT1(16'b0101010100000101),
    .MODE("LOGIC"))
    \_al_u2460|_al_u2525  (
    .a({_al_u2459_o,_al_u2524_o}),
    .b({open_n14581,\t/a/alu/n6 [6]}),
    .c({_al_u2126_o,_al_u2126_o}),
    .d({\t/a/alu/n6 [12],open_n14584}),
    .f({_al_u2460_o,_al_u2525_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    //.LUT1("~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .INIT_LUT0(16'b1010111110100000),
    .INIT_LUT1(16'b0001000111011101),
    .MODE("LOGIC"))
    \_al_u2462|_al_u2461  (
    .a({\t/a/alu/n35_lutinv ,\t/a/EX_A [13]}),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n14603}),
    .c({open_n14604,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n33_lutinv ,\t/a/EX_A [12]}),
    .f({_al_u2462_o,\t/a/alu/n35_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u2466|_al_u2464  (
    .a({_al_u2464_o,_al_u2372_o}),
    .b({\t/a/alu/n136_lutinv ,_al_u2463_o}),
    .c({_al_u2465_o,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }),
    .f({_al_u2466_o,_al_u2464_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*D*~A+C*~B*D*~A+~C*~B*D*A+C*~B*D*A"),
    //.LUTF1("0"),
    //.LUTG0("~C*~B*D*A+C*~B*D*A"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b0011001100000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0010001000000000),
    .INIT_LUTG1(16'b0011001100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2468|_al_u2488  (
    .a({\t/a/alu/n5 [11],\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .b({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .d({\t/a/EX_operation$0$_lutinv_placeOpt_3 ,_al_u2128_o}),
    .e({_al_u2128_o,\t/a/alu/n5 [9]}),
    .f({_al_u2468_o,_al_u2488_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUT1("(A*~(D*(B*~(C)*~(1)+~(B)*C*~(1)+B*C*~(1)+B*C*1)))"),
    .INIT_LUT0(16'b0001000011110000),
    .INIT_LUT1(16'b0010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2469 (
    .a({\t/a/EX_operation [1],\t/a/EX_A [11]}),
    .b({\t/a/EX_A [11],\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n14681,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .fx({open_n14686,_al_u2469_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*~A*D+C*~B*~A*D"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*~B*A*D+C*~B*A*D"),
    //.LUTG1("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0001000100010001),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0011001100110011),
    .INIT_LUTG1(16'b0101000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2470|_al_u2564  (
    .a({_al_u2469_o,_al_u2126_o}),
    .b({open_n14689,_al_u2563_o}),
    .c({\t/a/alu/n6 [11],open_n14690}),
    .e({_al_u2126_o,\t/a/alu/n6 [2]}),
    .f({_al_u2470_o,_al_u2564_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("~A*~D*~B*~C+A*~D*~B*~C+~A*~D*B*~C+A*~D*B*~C+~A*D*B*~C+A*D*B*~C+~A*~D*~B*C+A*~D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTG0("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG1("~A*~D*~B*~C+A*~D*~B*~C+~A*~D*~B*C+A*~D*~B*C"),
    .INIT_LUTF0(16'b1010101000000000),
    .INIT_LUTF1(16'b1100110011111111),
    .INIT_LUTG0(16'b1111111101010101),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2472|_al_u2471  (
    .a({open_n14715,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n14716}),
    .d({\t/a/alu/n36_lutinv ,\t/a/EX_A [12]}),
    .e({\t/a/alu/n34_lutinv ,\t/a/EX_A [11]}),
    .f({_al_u2472_o,\t/a/alu/n36_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u2476|_al_u2474  (
    .a({_al_u2474_o,_al_u2384_o}),
    .b({\t/a/alu/n135_lutinv ,_al_u2473_o}),
    .c({_al_u2475_o,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_1 }),
    .f({_al_u2476_o,_al_u2474_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUT1("(C*~(A*(D*~(B)*~(1)+~(D)*B*~(1)+D*B*~(1)+D*B*1)))"),
    .INIT_LUT0(16'b0001000011110000),
    .INIT_LUT1(16'b0111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2479 (
    .a({\t/a/EX_operation [2],\t/a/EX_A [10]}),
    .b({\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .d({\t/a/EX_A [10],\t/a/EX_operation [2]}),
    .mi({open_n14773,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .fx({open_n14778,_al_u2479_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+~A*C*~B*~D"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D"),
    //.LUTG0("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*~B*D+~A*C*~B*D"),
    //.LUTG1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D"),
    .INIT_LUTF0(16'b0000000000010001),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b0001000100010001),
    .INIT_LUTG1(16'b0011001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2480|_al_u2709  (
    .a({open_n14781,_al_u2708_o}),
    .b({_al_u2479_o,_al_u2479_o}),
    .d({_al_u2126_o,_al_u2126_o}),
    .e({\t/a/alu/n6 [10],\t/a/alu/n6 [10]}),
    .f({_al_u2480_o,_al_u2709_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*C*~B*~D+A*C*~B*~D+~A*C*B*~D+A*C*B*~D+~A*C*~B*D+A*C*~B*D+~A*C*B*D+A*C*B*D"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*~C*D+B*~A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG0("A*~C*~B*~D+A*C*~B*~D+A*~C*B*~D+A*C*B*~D+A*~C*~B*D+A*C*~B*D+A*~C*B*D+A*C*B*D"),
    //.LUTG1("~B*~A*~C*~D+B*~A*~C*~D+~B*~A*~C*D+B*~A*~C*D"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b1111010111110101),
    .INIT_LUTG0(16'b1010101010101010),
    .INIT_LUTG1(16'b0000010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2482|_al_u2481  (
    .a({\t/a/alu/n37_lutinv ,\t/a/EX_A [11]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [10]}),
    .e({\t/a/alu/n35_lutinv ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2482_o,\t/a/alu/n37_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*B*D+~A*C*B*D"),
    //.LUTF1("~A*~C*B*~D+~A*C*B*~D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG0("~A*~C*B*D+~A*C*B*D"),
    //.LUTG1("~A*~C*B*~D+~A*C*B*~D"),
    .INIT_LUTF0(16'b0100010011001100),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b0100010000000000),
    .INIT_LUTG1(16'b0000000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2486|_al_u2484  (
    .a({_al_u2484_o,_al_u2396_o}),
    .b({_al_u2485_o,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/alu/n134_lutinv ,_al_u2483_o}),
    .f({_al_u2486_o,_al_u2484_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*~C*D+~A*B*~C*D"),
    //.LUTG0("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0001000011110000),
    .INIT_LUTF1(16'b0000010100000101),
    .INIT_LUTG0(16'b0111000011110000),
    .INIT_LUTG1(16'b0101010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2490|_al_u2489  (
    .a({_al_u2489_o,\t/a/EX_A [9]}),
    .b({open_n14856,\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o }),
    .c({_al_u2126_o,\t/a/EX_operation [1]}),
    .d({open_n14859,\t/a/EX_operation [2]}),
    .e({\t/a/alu/n6 [9],\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .f({_al_u2490_o,_al_u2489_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    //.LUT1("~(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    .INIT_LUT0(16'b1100101011001010),
    .INIT_LUT1(16'b0101000001011111),
    .MODE("LOGIC"))
    \_al_u2492|_al_u2491  (
    .a({\t/a/alu/n36_lutinv ,\t/a/EX_A [9]}),
    .b({open_n14880,\t/a/EX_A [10]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n38_lutinv ,open_n14883}),
    .f({_al_u2492_o,\t/a/alu/n38_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*C*~A+B*~D*C*~A+~B*D*C*~A+B*D*C*~A+~B*~D*C*A+~B*D*C*A"),
    //.LUTF1("0"),
    //.LUTG0("~B*~D*C*A+~B*D*C*A"),
    //.LUTG1("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D"),
    .INIT_LUTF0(16'b0111000001110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0010000000100000),
    .INIT_LUTG1(16'b0000000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2496|_al_u2494  (
    .a({open_n14902,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 }),
    .b({_al_u2146_o,_al_u2409_o}),
    .c({\t/a/alu/n133_lutinv ,_al_u2161_o}),
    .d({_al_u2494_o,open_n14905}),
    .e({_al_u2495_o,_al_u2493_o}),
    .f({_al_u2496_o,_al_u2494_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    //.LUTG0("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    .INIT_LUTF0(16'b0001000011110000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b0111000011110000),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2500|_al_u2499  (
    .a({open_n14926,\t/a/EX_A [8]}),
    .b({_al_u2126_o,\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o }),
    .c({open_n14927,\t/a/EX_operation [1]}),
    .d({_al_u2499_o,\t/a/EX_operation [2]}),
    .e({\t/a/alu/n6 [8],\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .f({_al_u2500_o,_al_u2499_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)"),
    //.LUT1("~(A*~(D)*~(B)+A*D*~(B)+~(A)*D*B+A*D*B)"),
    .INIT_LUT0(16'b1110111001000100),
    .INIT_LUT1(16'b0001000111011101),
    .MODE("LOGIC"))
    \_al_u2502|_al_u2501  (
    .a({\t/a/alu/n39_lutinv ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [8]}),
    .d({\t/a/alu/n37_lutinv ,\t/a/EX_A [9]}),
    .f({_al_u2502_o,\t/a/alu/n39_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b1111101000001010),
    .MODE("LOGIC"))
    \_al_u2503|_al_u2544  (
    .a({_al_u2502_o,_al_u2502_o}),
    .b({open_n14972,_al_u2543_o}),
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_1 }),
    .d({_al_u2462_o,\t/a/EX_B [2]}),
    .f({_al_u2503_o,_al_u2544_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u2506|_al_u2504  (
    .a({_al_u2504_o,_al_u2421_o}),
    .b({\t/a/alu/n132_lutinv ,_al_u2503_o}),
    .c({_al_u2505_o,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2506_o,_al_u2504_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUT1("(B*~(D*(C*~(A)*~(1)+~(C)*A*~(1)+C*A*~(1)+C*A*1)))"),
    .INIT_LUT0(16'b0001000011110000),
    .INIT_LUT1(16'b0100110011001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2509 (
    .a({\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [7]}),
    .b({\t/a/EX_operation [1],\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_A [7],\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n15025,\t/a/EX_operation [0]}),
    .fx({open_n15030,_al_u2509_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*C*~B*~A+D*C*~B*~A+~D*C*B*~A+D*C*B*~A+~D*C*~B*A+D*C*~B*A+~D*C*B*A+D*C*B*A"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A"),
    //.LUTG0("~D*~C*~B*A+D*~C*~B*A+~D*C*~B*A+D*C*~B*A+~D*~C*B*A+D*~C*B*A+~D*C*B*A+D*C*B*A"),
    //.LUTG1("~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    .INIT_LUTF0(16'b1111000011110000),
    .INIT_LUTF1(16'b0101111101011111),
    .INIT_LUTG0(16'b1010101010101010),
    .INIT_LUTG1(16'b0101000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2512|_al_u2511  (
    .a({\t/a/alu/n38_lutinv ,\t/a/EX_A [8]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [7]}),
    .e({\t/a/alu/n40_lutinv ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2512_o,\t/a/alu/n40_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*~C*~A+D*B*~C*~A"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("~D*B*~C*~A+D*B*~C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D"),
    .INIT_LUTF0(16'b0000010000000100),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b0000111000001110),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2514|_al_u2513  (
    .a({open_n15059,\t/a/EX_B [2]}),
    .b({_al_u2161_o,_al_u2512_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_3 ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_3 }),
    .d({_al_u2513_o,open_n15062}),
    .e({_al_u2430_o,_al_u2472_o}),
    .f({_al_u2514_o,_al_u2513_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~C*A*~B+~D*C*A*~B+~D*~C*A*B+D*~C*A*B+~D*C*A*B+D*C*A*B"),
    //.LUTF1("A*~D*~B*~C+A*~D*B*~C+A*~D*~B*C+A*D*~B*C+A*~D*B*C+A*D*B*C"),
    //.LUTG0("D*~C*A*~B+D*C*A*~B+~D*~C*A*B+D*~C*A*B+~D*C*A*B+D*C*A*B"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b1010000010101010),
    .INIT_LUTG0(16'b1010101010001000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2516|_al_u2515  (
    .a({_al_u2515_o,_al_u2431_o}),
    .b({open_n15083,\t/a/EX_operation [0]}),
    .c({_al_u2334_o,open_n15084}),
    .d({_al_u2146_o,\t/a/EX_A [7]}),
    .e({_al_u2514_o,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2516_o,_al_u2515_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(A*~((~C*B))*~(0)+A*(~C*B)*~(0)+~(A)*(~C*B)*0+A*(~C*B)*0))"),
    //.LUT1("(~D*(A*~((~C*B))*~(1)+A*(~C*B)*~(1)+~(A)*(~C*B)*1+A*(~C*B)*1))"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2518 (
    .a({\t/a/alu/n5 [6],\t/a/alu/n5 [6]}),
    .b({\t/a/alu/n261_lutinv ,\t/a/alu/n261_lutinv }),
    .c({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .mi({open_n15119,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .fx({open_n15124,\t/a/alu/mux0_b6/B1_0 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+~A*B*C*~D+~A*B*~C*D+~A*B*C*D"),
    //.LUTF1("~C*~A*~B*~D+C*~A*~B*~D+~C*~A*B*~D+C*~A*B*~D+~C*A*B*~D+C*A*B*~D+~C*~A*~B*D+C*~A*~B*D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    //.LUTG0("A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~C*~A*~B*~D+C*~A*~B*~D+~C*~A*~B*D+C*~A*~B*D"),
    .INIT_LUTF0(16'b0100010001000100),
    .INIT_LUTF1(16'b1101110111011101),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0001000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2520|_al_u2519  (
    .a({\t/a/alu/n41_lutinv ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [6]}),
    .e({\t/a/alu/n39_lutinv ,\t/a/EX_A [7]}),
    .f({_al_u2520_o,\t/a/alu/n41_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*~A*~(0*B)))"),
    //.LUTF1("~B*~A*C*~D+~B*A*C*~D+B*~A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG0("(C*~(D*~A*~(1*B)))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1010000011110000),
    .INIT_LUTF1(16'b1111110000110000),
    .INIT_LUTG0(16'b1110000011110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2521|_al_u2523  (
    .a({open_n15153,_al_u2521_o}),
    .b({\t/a/EX_B [2],_al_u2443_o}),
    .c({_al_u2520_o,_al_u2522_o}),
    .d({_al_u2482_o,_al_u2161_o}),
    .e({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2521_o,_al_u2523_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(~(A)*~(B)*~(D)+~(A)*~(B)*D+A*~(B)*D+~(A)*B*D))"),
    //.LUT1("(D*~(~C*(B@A)))"),
    .INIT_LUT0(16'b0111000000010000),
    .INIT_LUT1(16'b1111100100000000),
    .MODE("LOGIC"))
    \_al_u2522|_al_u2526  (
    .a({\t/a/EX_A [6],\t/a/EX_A [6]}),
    .b({\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_operation [0],\t/a/EX_operation [1]}),
    .d({_al_u2431_o,\t/a/EX_operation [0]}),
    .f({_al_u2522_o,_al_u2526_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("(C*~(A*~D))"),
    //.LUTG0("0"),
    //.LUTG1("(C*~(A*~D))"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b1111000001010000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2524|_al_u2686  (
    .a({_al_u2146_o,_al_u2161_o}),
    .c({_al_u2523_o,open_n15198}),
    .d({_al_u2347_o,open_n15201}),
    .e({open_n15202,_al_u2187_o}),
    .f({_al_u2524_o,_al_u2686_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(A*~((~C*B))*~(0)+A*(~C*B)*~(0)+~(A)*(~C*B)*0+A*(~C*B)*0))"),
    //.LUT1("(~D*(A*~((~C*B))*~(1)+A*(~C*B)*~(1)+~(A)*(~C*B)*1+A*(~C*B)*1))"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2528 (
    .a({\t/a/alu/n5 [5],\t/a/alu/n5 [5]}),
    .b({\t/a/alu/n262_lutinv ,\t/a/alu/n262_lutinv }),
    .c({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .mi({open_n15235,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .fx({open_n15240,\t/a/alu/mux0_b5/B1_0 }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)"),
    //.LUT1("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT_LUT0(16'b1111101001010000),
    .INIT_LUT1(16'b0100011101000111),
    .MODE("LOGIC"))
    \_al_u2530|_al_u2529  (
    .a({\t/a/alu/n40_lutinv ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,open_n15243}),
    .c({\t/a/alu/n42_lutinv ,\t/a/EX_A [5]}),
    .d({open_n15246,\t/a/EX_A [6]}),
    .f({_al_u2530_o,\t/a/alu/n42_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u2532|_al_u2531  (
    .a({_al_u2531_o,_al_u2492_o}),
    .b({_al_u2453_o,_al_u2530_o}),
    .c({_al_u2161_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 }),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_2 ,\t/a/EX_B [2]}),
    .f({_al_u2532_o,_al_u2531_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(A*~(~C*(B@D)))"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1010100010100010),
    .MODE("LOGIC"))
    \_al_u2533|_al_u418  (
    .a({_al_u2431_o,\t/a/ID_rs1$0$_placeOpt_10 }),
    .b({\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ,\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/EX_operation [0],\t/a/regfile/regfile$4$ [5]}),
    .d({\t/a/EX_A [5],\t/a/regfile/regfile$5$ [5]}),
    .f({_al_u2533_o,_al_u418_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(D*~B))"),
    //.LUT1("(~A*~(C*~D))"),
    .INIT_LUT0(16'b0100000001010000),
    .INIT_LUT1(16'b0101010100000101),
    .MODE("LOGIC"))
    \_al_u2535|_al_u2534  (
    .a({_al_u2534_o,_al_u2532_o}),
    .b({open_n15305,_al_u2360_o}),
    .c({_al_u2126_o,_al_u2533_o}),
    .d({\t/a/alu/n6 [5],_al_u2146_o}),
    .f({_al_u2535_o,_al_u2534_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*A)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1010000010100000),
    .MODE("LOGIC"))
    \_al_u2538|_al_u2707  (
    .a({\t/a/alu/n263_lutinv ,open_n15326}),
    .c({_al_u2161_o,_al_u2161_o}),
    .d({open_n15331,_al_u2279_o}),
    .f({_al_u2538_o,_al_u2707_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*(~(A)*~(B)*~(0)+~(A)*~(B)*0+A*~(B)*0+~(A)*B*0)))"),
    //.LUT1("(A*~(C*(~(D)*~(B)*~(1)+~(D)*~(B)*1+D*~(B)*1+~(D)*B*1)))"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1000101000001010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2539 (
    .a({\t/a/EX_operation [2],\t/a/EX_A [4]}),
    .b({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .d({\t/a/EX_A [4],\t/a/EX_operation [2]}),
    .mi({open_n15362,\t/a/EX_operation [0]}),
    .fx({open_n15367,_al_u2539_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~D*~(~B*~(~0*A))))"),
    //.LUT1("(C*~(~D*~(~B*~(~1*A))))"),
    .INIT_LUT0(16'b1111000000010000),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2541 (
    .a({\t/a/alu/n5 [4],\t/a/alu/n5 [4]}),
    .b({_al_u2538_o,_al_u2538_o}),
    .c({_al_u2540_o,_al_u2540_o}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .mi({open_n15382,\t/a/EX_operation$0$_lutinv_placeOpt_2 }),
    .fx({open_n15387,_al_u2541_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C)"),
    //.LUT1("(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C)"),
    .INIT_LUT0(16'b1111101000001010),
    .INIT_LUT1(16'b1010111110100000),
    .MODE("LOGIC"))
    \_al_u2542|_al_u2550  (
    .a({\t/a/EX_A [5],\t/a/EX_A [3]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_A [4],\t/a/EX_A [4]}),
    .f({\t/a/alu/n43_lutinv ,\t/a/alu/n44_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*C*~D*~(A*~B))"),
    //.LUTF1("A*~B*~D*~C+A*~B*D*~C+A*~B*~D*C+A*~B*D*C"),
    //.LUTG0("(1*C*~D*~(A*~B))"),
    //.LUTG1("A*~B*~D*~C+A*~B*D*~C"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0010001000100010),
    .INIT_LUTG0(16'b0000000011010000),
    .INIT_LUTG1(16'b0000001000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2545|_al_u2547  (
    .a({_al_u2161_o,_al_u2146_o}),
    .b({_al_u2544_o,_al_u2373_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,_al_u2546_o}),
    .d({open_n15414,_al_u2545_o}),
    .e({_al_u2463_o,\t/a/EX_operation [2]}),
    .f({_al_u2545_o,_al_u2547_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*C)"),
    //.LUTF1("0"),
    //.LUTG0("(~B*C)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D"),
    .INIT_LUTF0(16'b0011000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0011000000110000),
    .INIT_LUTG1(16'b0000111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u254|_al_u1046  (
    .b({open_n15437,\t/a/WB_rd [0]}),
    .c({\t/a/WB_rd [4],\t/a/ID_rs2$0$_placeOpt_21 }),
    .e({\t/a/WB_regwritecs ,open_n15442}),
    .f({_al_u254_o,_al_u1046_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(0)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(0)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*0+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*0)"),
    //.LUTF1("~A*B*~D*~C+~A*B*D*~C+~A*B*~D*C+A*B*~D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(1)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(1)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*1+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*1)"),
    //.LUTG1("~A*B*~D*~C+~A*B*D*~C"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b1100010011000100),
    .INIT_LUTG0(16'b1010101010101010),
    .INIT_LUTG1(16'b0000010000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2552|_al_u2551  (
    .a({_al_u2551_o,_al_u2512_o}),
    .b({_al_u2161_o,\t/a/alu/n42_lutinv }),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_3 ,\t/a/alu/n44_lutinv }),
    .d({open_n15465,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({_al_u2473_o,\t/a/EX_B [2]}),
    .f({_al_u2552_o,_al_u2551_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~D*(C@A)))"),
    //.LUT1("(A*~B*~(D*~C))"),
    .INIT_LUT0(16'b1100110010000100),
    .INIT_LUT1(16'b0010000000100010),
    .MODE("LOGIC"))
    \_al_u2554|_al_u2553  (
    .a({_al_u2553_o,\t/a/EX_A [3]}),
    .b({_al_u2552_o,_al_u2431_o}),
    .c({_al_u2385_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_1 }),
    .d({_al_u2146_o,\t/a/EX_operation [0]}),
    .f({_al_u2554_o,_al_u2553_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(0)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(0)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*0+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*0)"),
    //.LUT1("(~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(A)*~(1)+~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A*~(1)+~(~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*A*1+~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*A*1)"),
    .INIT_LUT0(16'b0011001100001111),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2560 (
    .a({_al_u2520_o,_al_u2520_o}),
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/alu/n43_lutinv }),
    .c({\t/a/alu/n45_lutinv ,\t/a/alu/n45_lutinv }),
    .d({\t/a/alu/n43_lutinv ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .mi({open_n15518,\t/a/EX_B [2]}),
    .fx({open_n15523,_al_u2560_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~A*B*~D+C*~A*B*~D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    //.LUTF1("~B*~C*~D*A+B*~C*~D*A+~B*C*~D*A+B*C*~D*A+B*~C*D*A+B*C*D*A"),
    //.LUTG0("~C*~A*B*D+C*~A*B*D"),
    //.LUTG1("B*~C*~D*A+B*C*~D*A+~B*~C*D*A+B*~C*D*A+~B*C*D*A+B*C*D*A"),
    .INIT_LUTF0(16'b1100110001000100),
    .INIT_LUTF1(16'b1000100010101010),
    .INIT_LUTG0(16'b0100010000000000),
    .INIT_LUTG1(16'b1010101010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2561|_al_u2565  (
    .a({_al_u2431_o,\t/a/EX_B [2]}),
    .b({\t/a/EX_operation [0],\t/a/EX_operation [1]}),
    .d({\t/a/EX_B [2],\t/a/EX_operation [0]}),
    .e({\t/a/EX_A [2],\t/a/EX_A [2]}),
    .f({_al_u2561_o,_al_u2565_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*~(B*~(A)*~(0)+B*A*~(0)+~(B)*A*0+B*A*0)))"),
    //.LUTF1("(D*~(B*~C))"),
    //.LUTG0("(C*~(D*~(B*~(A)*~(1)+B*A*~(1)+~(B)*A*1+B*A*1)))"),
    //.LUTG1("(D*~(B*~C))"),
    .INIT_LUTF0(16'b1100000011110000),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b1010000011110000),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2563|_al_u2562  (
    .a({open_n15550,_al_u2483_o}),
    .b({_al_u2146_o,_al_u2560_o}),
    .c({_al_u2397_o,_al_u2561_o}),
    .d({_al_u2562_o,_al_u2161_o}),
    .e({open_n15553,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2563_o,_al_u2562_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*B*A)"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D"),
    //.LUTG0("(~1*~D*~C*B*A)"),
    //.LUTG1("~A*~B*C*~D+~A*B*C*~D"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2568|_al_u2567  (
    .a({_al_u2567_o,_al_u2184_o}),
    .b({open_n15574,_al_u2161_o}),
    .c({\t/a/EX_operation$0$_lutinv_placeOpt_2 ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_operation [1],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/alu/n5 [0],\t/a/EX_B [2]}),
    .f({_al_u2568_o,_al_u2567_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*(~(A)*~(B)*~(0)+~(A)*~(B)*0+A*~(B)*0+~(A)*B*0))"),
    //.LUT1("(D*C*(~(B)*~(A)*~(1)+~(B)*~(A)*1+B*~(A)*1+~(B)*A*1))"),
    .INIT_LUT0(16'b0001000000000000),
    .INIT_LUT1(16'b0111000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2569 (
    .a({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [0]}),
    .b({\t/a/EX_A [0],\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n15609,\t/a/EX_operation [0]}),
    .fx({open_n15614,_al_u2569_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+A*B*~C*~D+~A*B*~C*D+A*B*~C*D"),
    //.LUTF1("(A*C)"),
    //.LUTG0("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG1("(A*C)"),
    .INIT_LUTF0(16'b0000110000001100),
    .INIT_LUTF1(16'b1010000010100000),
    .INIT_LUTG0(16'b0000000011001100),
    .INIT_LUTG1(16'b1010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u256|_al_u1712  (
    .a({\t/a/WB_regwritecs ,open_n15617}),
    .b({open_n15618,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/WB_rd [4],\t/a/regfile/regfile$22$ [0]}),
    .d({open_n15621,\t/a/regfile/regfile$23$ [0]}),
    .e({open_n15622,\t/a/ID_rs2$0$_placeOpt_21 }),
    .f({_al_u256_o,_al_u1712_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+~A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTF1("(~C*~(~0*~(~B*~(D*~A))))"),
    //.LUTG0("0"),
    //.LUTG1("(~C*~(~1*~(~B*~(D*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100010001),
    .INIT_LUTF1(16'b0000001000000011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2570|t/a/ex_mem/reg4_b0  (
    .a({\t/a/alu/n8 ,_al_u2128_o}),
    .b({_al_u2568_o,_al_u2571_o}),
    .c({_al_u2569_o,open_n15643}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [1],_al_u2570_o}),
    .e({\t/a/EX_operation [2],_al_u2577_o}),
    .sr(rst_pad),
    .f({_al_u2570_o,\t/a/aludat [0]}),
    .q({open_n15662,\t/a/MEM_aludat [0]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(B*~D))"),
    //.LUTF1("(A*~B)"),
    //.LUTG0("(~A*~(B*~D))"),
    //.LUTG1("(A*~B)"),
    .INIT_LUTF0(16'b0101010100010001),
    .INIT_LUTF1(16'b0010001000100010),
    .INIT_LUTG0(16'b0101010100010001),
    .INIT_LUTG1(16'b0010001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2571|_al_u2510  (
    .a({_al_u2126_o,_al_u2509_o}),
    .b({\t/a/alu/n6 [0],_al_u2126_o}),
    .d({open_n15667,\t/a/alu/n6 [7]}),
    .f({_al_u2571_o,_al_u2510_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+~A*C*B*D"),
    //.LUTF1("0"),
    //.LUTG0("~A*~C*B*~D+~A*C*B*~D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    .INIT_LUTF0(16'b0111011101110111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0100010001000100),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2572|_al_u2543  (
    .a({open_n15690,\t/a/alu/n41_lutinv }),
    .b({open_n15691,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2543_o,open_n15696}),
    .e({\t/a/EX_B [2],\t/a/alu/n43_lutinv }),
    .f({_al_u2572_o,_al_u2543_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(A*C)"),
    //.LUTG0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("(A*C)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010000010100000),
    .INIT_LUTG0(16'b0101010101010101),
    .INIT_LUTG1(16'b1010000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2573|_al_u2184  (
    .a({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_A [1],open_n15719}),
    .e({open_n15724,\t/a/EX_A [0]}),
    .f({_al_u2573_o,_al_u2184_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D))"),
    //.LUTF1("(A*~((~D*~B)*~(C)*~(0)+(~D*~B)*C*~(0)+~((~D*~B))*C*0+(~D*~B)*C*0))"),
    //.LUTG0("(~1*(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D))"),
    //.LUTG1("(A*~((~D*~B)*~(C)*~(1)+(~D*~B)*C*~(1)+~((~D*~B))*C*1+(~D*~B)*C*1))"),
    .INIT_LUTF0(16'b1010101011111100),
    .INIT_LUTF1(16'b1010101010001000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2575|_al_u2574  (
    .a({_al_u2161_o,\t/a/alu/n45_lutinv }),
    .b({_al_u2572_o,_al_u2573_o}),
    .c({_al_u2503_o,_al_u2184_o}),
    .d({_al_u2574_o,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_1 ,\t/a/EX_B [2]}),
    .f({_al_u2575_o,_al_u2574_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~D*(C@A)))"),
    //.LUT1("(A*~B*~(D*~C))"),
    .INIT_LUT0(16'b1100110010000100),
    .INIT_LUT1(16'b0010000000100010),
    .MODE("LOGIC"))
    \_al_u2577|_al_u2576  (
    .a({_al_u2576_o,\t/a/EX_A [0]}),
    .b({_al_u2575_o,_al_u2431_o}),
    .c({_al_u2422_o,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2146_o,\t/a/EX_operation$0$_lutinv_placeOpt_2 }),
    .f({_al_u2577_o,_al_u2576_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0011001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2580|_al_u2230  (
    .b({_al_u2530_o,open_n15789}),
    .c({open_n15790,\t/a/EX_B [2]}),
    .d({open_n15793,_al_u2229_o}),
    .e({\t/a/EX_B [2],open_n15794}),
    .f({_al_u2580_o,\t/a/alu/n105_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000010100000011),
    .INIT_LUTF1(16'b0000000011001111),
    .INIT_LUTG0(16'b0000010100000011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2582|_al_u2581  (
    .a({open_n15815,\t/a/EX_A [2]}),
    .b({\t/a/alu/n44_lutinv ,\t/a/EX_A [1]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2581_o,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/EX_B [2],open_n15818}),
    .f({_al_u2582_o,_al_u2581_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~((~C*~B)*~(A)*~(0)+(~C*~B)*A*~(0)+~((~C*~B))*A*0+(~C*~B)*A*0))"),
    //.LUT1("(D*~((~C*~B)*~(A)*~(1)+(~C*~B)*A*~(1)+~((~C*~B))*A*1+(~C*~B)*A*1))"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b0101010100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2583 (
    .a({_al_u2493_o,_al_u2493_o}),
    .b({_al_u2580_o,_al_u2580_o}),
    .c({_al_u2582_o,_al_u2582_o}),
    .d({_al_u2161_o,_al_u2161_o}),
    .mi({open_n15851,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_3 }),
    .fx({open_n15856,_al_u2583_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+A*~B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~C*~B*~D*A+C*~B*~D*A+~C*B*~D*A+C*B*~D*A+~C*B*D*A+C*B*D*A"),
    //.LUTG0("~A*~B*C*D+A*~B*C*D"),
    //.LUTG1("~C*B*~D*A+C*B*~D*A+~C*~B*D*A+C*~B*D*A+~C*B*D*A+C*B*D*A"),
    .INIT_LUTF0(16'b1111000000110000),
    .INIT_LUTF1(16'b1000100010101010),
    .INIT_LUTG0(16'b0011000000000000),
    .INIT_LUTG1(16'b1010101010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2584|_al_u2587  (
    .a({_al_u2431_o,open_n15859}),
    .b({\t/a/EX_operation [0],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .c({open_n15860,\t/a/EX_operation [1]}),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation [0]}),
    .e({\t/a/EX_A [1],\t/a/EX_A [1]}),
    .f({_al_u2584_o,_al_u2587_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("C*~B*~D*~A+C*~B*D*~A"),
    //.LUTG0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("C*~B*~D*~A+C*~B*D*~A+C*~B*~D*A+C*~B*D*A"),
    .INIT_LUTF0(16'b0101010001010100),
    .INIT_LUTF1(16'b0001000000010000),
    .INIT_LUTG0(16'b0101010101010101),
    .INIT_LUTG1(16'b0011000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2585|_al_u2586  (
    .a({_al_u2146_o,_al_u2585_o}),
    .b({_al_u2583_o,\t/a/alu/n6 [1]}),
    .c({_al_u2584_o,_al_u2128_o}),
    .e({_al_u2410_o,\t/a/EX_operation$0$_lutinv_placeOpt_3 }),
    .f({_al_u2585_o,_al_u2586_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUT1("(A*~(~D*~(~C*~B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111001001010000),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2589|t/a/mem_wb/reg0_b6  (
    .a({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({i_data[3],_al_u1908_o}),
    .c({i_data[6],\t/a/MEM_aludat [6]}),
    .clk(clock_pad),
    .d({_al_u1908_o,i_data[6]}),
    .sr(rst_pad),
    .f({_al_u2589_o,open_n15920}),
    .q({open_n15924,\t/a/reg_writedat [6]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUT1("(~A*~(~D*~C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111001001010000),
    .INIT_LUT1(16'b0101010101010100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2590|t/a/mem_wb/reg0_b5  (
    .a({_al_u1908_o,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({i_data[0],_al_u1908_o}),
    .c({i_data[5],\t/a/MEM_aludat [5]}),
    .clk(clock_pad),
    .d({i_data[4],i_data[5]}),
    .sr(rst_pad),
    .f({_al_u2590_o,open_n15938}),
    .q({open_n15942,\t/a/reg_writedat [5]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*~B*~(~0*A))"),
    //.LUT1("(~D*C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000000010000),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2591 (
    .a({\t/a/mux4_b7/B0_0 ,\t/a/mux4_b7/B0_0 }),
    .b({_al_u1904_o,_al_u1904_o}),
    .c({_al_u2589_o,_al_u2589_o}),
    .d({_al_u2590_o,_al_u2590_o}),
    .mi({open_n15955,_al_u1908_o}),
    .fx({open_n15960,_al_u2591_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~0*~D*~C*~B))"),
    //.LUT1("(C*~(~1*~D*~A*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101010101000),
    .INIT_LUT1(16'b1111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    _al_u2592 (
    .a({i_data[31],_al_u1918_o}),
    .b({i_data[27],i_data[27]}),
    .c({_al_u1918_o,i_data[31]}),
    .clk(clock_pad),
    .d({i_data[29],i_data[29]}),
    .mi(i_data[29:28]),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .fx({open_n15977,_al_u2592_o}),
    .q({\trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/level_0_r ,open_n15978}));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~A*B*~D+C*~A*B*~D+~C*A*B*~D+C*A*B*~D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    //.LUTF1("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D+~C*B*A*~D+C*B*A*~D+~C*B*~A*D+C*B*~A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG0("~C*~A*~B*D+C*~A*~B*D+~C*~A*B*D+C*~A*B*D"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110011001100),
    .INIT_LUTF1(16'b1100110011011101),
    .INIT_LUTG0(16'b0101010100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2593|t/a/mem_wb/reg0_b1  (
    .a({i_data[2],_al_u1908_o}),
    .b({_al_u1908_o,\t/a/MEM_aludat [1]}),
    .clk(clock_pad),
    .d({i_data[1],i_data[1]}),
    .e({_al_u1940_o,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .sr(rst_pad),
    .f({_al_u2593_o,open_n15996}),
    .q({open_n16000,\t/a/reg_writedat [1]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*~C))"),
    //.LUT1("(~B*C*~D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111111101110),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2594|t/a/mem_wb/reg0_b8  (
    .a({_al_u2591_o,_al_u1902_o}),
    .b({_al_u1906_o,_al_u1906_o}),
    .c({_al_u2593_o,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({_al_u2592_o,\t/a/MEM_aludat [8]}),
    .sr(rst_pad),
    .f({_al_u2594_o,open_n16014}),
    .q({open_n16018,\t/a/reg_writedat [8]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("(~B*~(~A*~C))"),
    //.LUTG0("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("(~B*~(~A*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0011001000110010),
    .INIT_LUTG0(16'b1111000011110000),
    .INIT_LUTG1(16'b0011001000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2595|_al_u2890  (
    .a({i_data[13],\t/a/instr/n12 [0]}),
    .b({_al_u1903_o,open_n16019}),
    .c({i_data[14],\t/memstraddress [0]}),
    .clk(clock_pad),
    .e({open_n16023,_al_u2109_o}),
    .mi({i_data[14],i_data[14]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u2595_o,_al_u2890_o}),
    .q({\trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*~(~C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100010101000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2597|_al_u1964  (
    .a({_al_u1918_o,_al_u1950_o}),
    .b({i_data[26],\t/busarbitration/n3_placeOpt_2 }),
    .c({i_data[30],\t/busarbitration/instruction [30]}),
    .clk(clock_pad),
    .d({open_n16040,i_data[30]}),
    .mi({i_data[30],i_data[30]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({_al_u2597_o,\t/a/IF_skip_addr [10]}),
    .q({\trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~0*~D*~C*~B))"),
    //.LUT1("(A*~(~1*~D*~C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101010101000),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    _al_u2598 (
    .a({_al_u1918_o,_al_u1918_o}),
    .b({i_data[18],i_data[18]}),
    .c({i_data[16],i_data[16]}),
    .clk(clock_pad),
    .d({i_data[23],i_data[23]}),
    .mi({i_data[23],i_data[21]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .fx({open_n16068,_al_u2598_o}),
    .q({\trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/level_0_r ,open_n16069}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*A)"),
    //.LUT1("(~1*~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2599 (
    .a({_al_u2594_o,_al_u2594_o}),
    .b({_al_u2595_o,_al_u2595_o}),
    .c({_al_u2596_o,_al_u2596_o}),
    .d({_al_u2597_o,_al_u2597_o}),
    .mi({open_n16082,_al_u2598_o}),
    .fx({open_n16087,_al_u2599_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    //.LUT1("(D*~(~B*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101010011),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2600|_al_u1962  (
    .a({open_n16090,i_data[20]}),
    .b({i_data[20],\t/busarbitration/instruction [20]}),
    .c({i_data[22],\t/busarbitration/n3_placeOpt_5 }),
    .clk(clock_pad),
    .d({_al_u1918_o,open_n16092}),
    .mi({i_data[22],i_data[22]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u2600_o,_al_u1962_o}),
    .q({\trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D*A)"),
    //.LUTF1("(~C*~A*~(B*~(~0*~D)))"),
    //.LUTG0("(C*D*A)"),
    //.LUTG1("(~C*~A*~(B*~(~1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010000000000000),
    .INIT_LUTF1(16'b0000000100000101),
    .INIT_LUTG0(16'b1010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2601|t/a/instr/instr_nop_reg  (
    .a({_al_u2600_o,_al_u2599_o}),
    .b({_al_u1918_o,open_n16106}),
    .c({_al_u1917_o,_al_u2602_o}),
    .clk(clock_pad),
    .d({i_data[25],_al_u2601_o}),
    .e({i_data[24],open_n16108}),
    .sr(rst_pad),
    .f({_al_u2601_o,open_n16123}),
    .q({open_n16127,\t/instrnop }));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*~C))"),
    //.LUT1("(~B*~(A*~(~D*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111111101110),
    .INIT_LUT1(16'b0001000100010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2602|t/a/mem_wb/reg0_b15  (
    .a({_al_u1918_o,_al_u1917_o}),
    .b({_al_u1935_o,_al_u1935_o}),
    .c({i_data[19],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({i_data[17],\t/a/MEM_aludat [15]}),
    .sr(rst_pad),
    .f({_al_u2602_o,open_n16141}),
    .q({open_n16145,\t/a/reg_writedat [15]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(B*A)"),
    //.LUTG0("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("(B*A)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1000100010001000),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2605|_al_u1799  (
    .a({_al_u1797_o,open_n16146}),
    .b({\t/a/condition/n1_lutinv ,_al_u1798_o}),
    .e({open_n16153,\t/a/n9_lutinv }),
    .f({\t/a/risk_jump/n19 ,\t/a/alu_A_select [0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~0*~D*C*B))"),
    //.LUT1("(~B*~(~1*~C*D*A))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0011001100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2606 (
    .a({\t/a/risk_jump/n19 ,_al_u2604_o}),
    .b({_al_u2604_o,\t/a/risk_jump/n19 }),
    .c({\t/a/risk_jump/n35_lutinv ,\t/a/risk_jump/n42_lutinv }),
    .d({\t/a/risk_jump/n42_lutinv ,\t/a/risk_jump/n35_lutinv }),
    .mi({open_n16186,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .fx({open_n16191,_al_u2606_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~0*~D*C*B))"),
    //.LUT1("(~A*~(~1*~D*C*B))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0101010101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2606_placeOpt_1 (
    .a({_al_u2604_o,_al_u2604_o}),
    .b({\t/a/risk_jump/n19 ,\t/a/risk_jump/n19 }),
    .c({\t/a/risk_jump/n42_lutinv ,\t/a/risk_jump/n42_lutinv }),
    .d({\t/a/risk_jump/n35_lutinv ,\t/a/risk_jump/n35_lutinv }),
    .mi({open_n16206,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .fx({open_n16211,_al_u2606_o_placeOpt_1}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~0*~D*C*B))"),
    //.LUT1("(~A*~(~1*~D*C*B))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0101010101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2606_placeOpt_2 (
    .a({_al_u2604_o,_al_u2604_o}),
    .b({\t/a/risk_jump/n19 ,\t/a/risk_jump/n19 }),
    .c({\t/a/risk_jump/n42_lutinv ,\t/a/risk_jump/n42_lutinv }),
    .d({\t/a/risk_jump/n35_lutinv ,\t/a/risk_jump/n35_lutinv }),
    .mi({open_n16226,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .fx({open_n16231,_al_u2606_o_placeOpt_2}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~0*~D*C*B))"),
    //.LUT1("(~A*~(~1*~D*C*B))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0101010101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2606_placeOpt_3 (
    .a({_al_u2604_o,_al_u2604_o}),
    .b({\t/a/risk_jump/n19 ,\t/a/risk_jump/n19 }),
    .c({\t/a/risk_jump/n42_lutinv ,\t/a/risk_jump/n42_lutinv }),
    .d({\t/a/risk_jump/n35_lutinv ,\t/a/risk_jump/n35_lutinv }),
    .mi({open_n16246,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .fx({open_n16251,_al_u2606_o_placeOpt_3}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*~A)"),
    //.LUTF1("(~D*~C)"),
    //.LUTG0("(~1*~D*~C*~B*~A)"),
    //.LUTG1("(~D*~C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2608|t/a/ex_mem/reg0_b0  (
    .a({open_n16254,\t/a/EX_rd [0]}),
    .b({open_n16255,\t/a/EX_rd [1]}),
    .c({\t/a/aluin/n11_lutinv ,\t/a/EX_rd [2]}),
    .clk(clock_pad),
    .d({_al_u2607_o,\t/a/EX_rd [3]}),
    .e({open_n16257,\t/a/EX_rd [4]}),
    .mi({open_n16259,\t/a/EX_rd [0]}),
    .sr(rst_pad),
    .f({_al_u2608_o,_al_u2607_o}),
    .q({open_n16274,\t/a/MEM_rd [0]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(~B*~C)"),
    //.LUTG0("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG1("(~B*~C)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000001100000011),
    .INIT_LUTG0(16'b1101110111011101),
    .INIT_LUTG1(16'b0000001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2610|_al_u2710  (
    .a({open_n16275,_al_u2610_o_placeOpt_1}),
    .b({_al_u2604_o,\t/a/ID_read_dat2 [10]}),
    .c({_al_u2609_o,open_n16276}),
    .e({open_n16281,_al_u2606_o_placeOpt_1}),
    .f({_al_u2610_o,_al_u2710_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("(~C*~A)"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("(~C*~A)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000010100000101),
    .INIT_LUTG0(16'b1111001111110011),
    .INIT_LUTG1(16'b0000010100000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2610|_al_u2710_placeOpt_1  (
    .a({_al_u2609_o,open_n16302}),
    .b({open_n16303,_al_u2610_o}),
    .c({_al_u2604_o,\t/a/ID_read_dat2 [10]}),
    .e({open_n16308,_al_u2606_o_placeOpt_1}),
    .f({_al_u2610_o_placeOpt_1,open_n16324}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTF1("(~A*~D)"),
    //.LUTG0("~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG1("(~A*~D)"),
    .INIT_LUTF0(16'b1010101010101010),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b1010000010100000),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2610|_al_u2710_placeOpt_2  (
    .a({_al_u2604_o,_al_u2606_o_placeOpt_1}),
    .c({open_n16332,\t/a/ID_read_dat2 [10]}),
    .d({_al_u2609_o,open_n16335}),
    .e({open_n16336,_al_u2610_o_placeOpt_1}),
    .f({_al_u2610_o_placeOpt_2,open_n16352}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~A*B))"),
    //.LUTF1("(~A*~D)"),
    //.LUTG0("(D*~(~A*B))"),
    //.LUTG1("(~A*~D)"),
    .INIT_LUTF0(16'b1011101100000000),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b1011101100000000),
    .INIT_LUTG1(16'b0000000001010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2610|_al_u2710_placeOpt_3  (
    .a({_al_u2604_o,\t/a/ID_read_dat2 [10]}),
    .b({open_n16358,_al_u2610_o_placeOpt_1}),
    .d({_al_u2609_o,_al_u2606_o_placeOpt_1}),
    .f({_al_u2610_o_placeOpt_3,open_n16380}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~A*~(C*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~A*~(C*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1010101011101010),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111101011101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2612|t/a/regfile/reg0_b127  (
    .a({_al_u2611_o,_al_u2606_o_placeOpt_1}),
    .b({\t/a/aludat [31],_al_u2610_o_placeOpt_1}),
    .c({_al_u2606_o_placeOpt_1,\t/a/MEM_aludat [31]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o_placeOpt_1,\t/a/reg_writedat [31]}),
    .e({\t/a/ID_read_dat2 [31],open_n16386}),
    .mi({open_n16388,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [31],_al_u2611_o}),
    .q({open_n16403,\t/a/regfile/regfile$3$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~0*~D*C*B))"),
    //.LUT1("(~A*~(~1*~C*D*B))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0101010101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2614 (
    .a({_al_u2613_o,_al_u2613_o}),
    .b({\t/a/risk_jump/n19 ,\t/a/risk_jump/n19 }),
    .c({\t/a/risk_jump/n11_lutinv ,\t/a/risk_jump/n24_lutinv }),
    .d({\t/a/risk_jump/n24_lutinv ,\t/a/risk_jump/n11_lutinv }),
    .mi({open_n16416,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .fx({open_n16421,_al_u2614_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~0*~D*C*B))"),
    //.LUT1("(~A*~(~1*~C*D*B))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0101010101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2614_placeOpt_1 (
    .a({_al_u2613_o,_al_u2613_o}),
    .b({\t/a/risk_jump/n19 ,\t/a/risk_jump/n19 }),
    .c({\t/a/risk_jump/n11_lutinv ,\t/a/risk_jump/n24_lutinv }),
    .d({\t/a/risk_jump/n24_lutinv ,\t/a/risk_jump/n11_lutinv }),
    .mi({open_n16436,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .fx({open_n16441,_al_u2614_o_placeOpt_1}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~0*~D*C*B))"),
    //.LUT1("(~B*~(~1*~D*C*A))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0011001100110011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2614_placeOpt_2 (
    .a({\t/a/risk_jump/n19 ,_al_u2613_o}),
    .b({_al_u2613_o,\t/a/risk_jump/n19 }),
    .c({\t/a/risk_jump/n24_lutinv ,\t/a/risk_jump/n24_lutinv }),
    .d({\t/a/risk_jump/n11_lutinv ,\t/a/risk_jump/n11_lutinv }),
    .mi({open_n16456,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .fx({open_n16461,_al_u2614_o_placeOpt_2}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~0*~D*C*B))"),
    //.LUT1("(~A*~(~1*~C*D*B))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0101010101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2614_placeOpt_3 (
    .a({_al_u2613_o,_al_u2613_o}),
    .b({\t/a/risk_jump/n19 ,\t/a/risk_jump/n19 }),
    .c({\t/a/risk_jump/n11_lutinv ,\t/a/risk_jump/n24_lutinv }),
    .d({\t/a/risk_jump/n24_lutinv ,\t/a/risk_jump/n11_lutinv }),
    .mi({open_n16476,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .fx({open_n16481,_al_u2614_o_placeOpt_3}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~B*A))"),
    //.LUTF1("(~D*~B)"),
    //.LUTG0("(D*~(~B*A))"),
    //.LUTG1("(~D*~B)"),
    .INIT_LUTF0(16'b1101110100000000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b1101110100000000),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2616|_al_u2692  (
    .a({open_n16484,_al_u2616_o}),
    .b({_al_u2615_o,\t/a/ID_read_dat1 [14]}),
    .d({_al_u2613_o,_al_u2614_o_placeOpt_1}),
    .f({_al_u2616_o,_al_u2692_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0010001000100010),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b1010101010101010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2616|_al_u2692_placeOpt_1  (
    .a({open_n16511,_al_u2614_o_placeOpt_1}),
    .b({open_n16512,_al_u2616_o}),
    .d({_al_u2613_o,open_n16517}),
    .e({_al_u2615_o,\t/a/ID_read_dat1 [14]}),
    .f({_al_u2616_o_placeOpt_1,open_n16533}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0011001100000000),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2616|_al_u2692_placeOpt_2  (
    .a({_al_u2615_o,open_n16539}),
    .b({open_n16540,_al_u2616_o}),
    .d({open_n16545,_al_u2614_o_placeOpt_1}),
    .e({_al_u2613_o,\t/a/ID_read_dat1 [14]}),
    .f({_al_u2616_o_placeOpt_2,open_n16561}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0011001100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2616|_al_u2692_placeOpt_3  (
    .b({open_n16569,_al_u2616_o}),
    .c({_al_u2613_o,open_n16570}),
    .d({_al_u2615_o,_al_u2614_o_placeOpt_1}),
    .e({open_n16573,\t/a/ID_read_dat1 [14]}),
    .f({_al_u2616_o_placeOpt_3,open_n16589}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*~C*~D+~B*A*~C*~D+~B*~A*~C*D+B*~A*~C*D+~B*A*~C*D+B*A*~C*D+B*~A*C*D+B*A*C*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("B*~A*~C*D+B*A*~C*D+B*~A*C*D+B*A*C*D"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b1110110011101100),
    .INIT_LUTG0(16'b1100110000000000),
    .INIT_LUTG1(16'b1111110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2618|t/a/id_ex/reg8_b31  (
    .a({\t/a/aludat [31],open_n16595}),
    .b({_al_u2617_o,_al_u333_o}),
    .c({_al_u2614_o_placeOpt_1,_al_u500_o}),
    .clk(clock_pad),
    .d({\t/a/ID_read_dat1 [31],\t/a/reg_writedat [31]}),
    .e({_al_u2616_o_placeOpt_2,_al_u490_o}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [31],\t/a/ID_read_dat1 [31]}),
    .q({open_n16614,\t/a/EX_regdat1 [31]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(A*(C*~(1)*~(D)+C*1*~(D)+~(C)*1*D+C*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1110111011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2622 (
    .a({_al_u2614_o_placeOpt_2,\t/a/aludat [30]}),
    .b({_al_u2621_o,_al_u2621_o}),
    .c({\t/a/aludat [30],_al_u2614_o_placeOpt_2}),
    .d({_al_u2616_o_placeOpt_2,_al_u2616_o_placeOpt_2}),
    .mi({open_n16627,\t/a/ID_read_dat1 [30]}),
    .fx({open_n16632,\t/a/ID_jump_regdat1 [30]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*~C*~D+~B*A*~C*~D+~B*~A*~C*D+B*~A*~C*D+~B*A*~C*D+B*A*~C*D+B*~A*C*D+B*A*C*D"),
    //.LUTF1("~A*B*C*~D+A*B*C*~D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("B*~A*~C*D+B*A*~C*D+B*~A*C*D+B*A*C*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b1010000011000000),
    .INIT_LUTG0(16'b1100110000000000),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2626|t/a/id_ex/reg8_b29  (
    .a({\t/a/ID_read_dat1 [29],open_n16635}),
    .b({\t/a/aludat [29],_al_u333_o}),
    .c({_al_u2614_o_placeOpt_2,_al_u563_o}),
    .clk(clock_pad),
    .d({_al_u2616_o_placeOpt_2,\t/a/reg_writedat [29]}),
    .e({_al_u2625_o,_al_u553_o}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [29],\t/a/ID_read_dat1 [29]}),
    .q({open_n16654,\t/a/EX_regdat1 [29]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~C*~A*D+~B*C*~A*D+~B*~C*A*D+~B*C*A*D"),
    //.LUTF1("~(~D*~(C*(A*~(0)*~(B)+A*0*~(B)+~(A)*0*B+A*0*B)))"),
    //.LUTG0("~B*~C*A*~D+~B*C*A*~D+~B*~C*A*D+~B*C*A*D"),
    //.LUTG1("~(~D*~(C*(A*~(1)*~(B)+A*1*~(B)+~(A)*1*B+A*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100000000),
    .INIT_LUTF1(16'b1111111100100000),
    .INIT_LUTG0(16'b0010001000100010),
    .INIT_LUTG1(16'b1111111111100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2628|t/a/regfile/reg0_b124  (
    .a({\t/a/aludat [28],\t/a/MEM_aludat [28]}),
    .b({_al_u2610_o_placeOpt_3,_al_u2606_o_placeOpt_3}),
    .c({_al_u2606_o_placeOpt_3,open_n16655}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2627_o,\t/a/reg_writedat [28]}),
    .e({\t/a/ID_read_dat2 [28],_al_u2610_o_placeOpt_3}),
    .mi({open_n16657,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [28],_al_u2627_o}),
    .q({open_n16672,\t/a/regfile/regfile$3$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+A*~C*B*D+A*C*B*D"),
    //.LUTF1("~A*B*C*~D+A*B*C*~D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("A*~C*~B*D+A*C*~B*D+A*~C*B*D+A*C*B*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101100010001),
    .INIT_LUTF1(16'b1010000011000000),
    .INIT_LUTG0(16'b1010101000000000),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2630|t/a/id_ex/reg8_b28  (
    .a({\t/a/ID_read_dat1 [28],_al_u333_o}),
    .b({\t/a/aludat [28],_al_u584_o}),
    .c({_al_u2614_o_placeOpt_2,open_n16673}),
    .clk(clock_pad),
    .d({_al_u2616_o_placeOpt_1,\t/a/reg_writedat [28]}),
    .e({_al_u2629_o,_al_u574_o}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [28],\t/a/ID_read_dat1 [28]}),
    .q({open_n16692,\t/a/EX_regdat1 [28]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*~A*C+~B*D*~A*C+~B*~D*A*C+~B*D*A*C"),
    //.LUTF1("~(~A*~(C*(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("~B*~D*A*~C+~B*D*A*~C+~B*~D*A*C+~B*D*A*C"),
    //.LUTG1("~(~A*~(C*(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000000110000),
    .INIT_LUTF1(16'b1011101010101010),
    .INIT_LUTG0(16'b0010001000100010),
    .INIT_LUTG1(16'b1111101011101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2632|t/a/regfile/reg0_b123  (
    .a({_al_u2631_o,\t/a/MEM_aludat [27]}),
    .b({_al_u2610_o_placeOpt_3,_al_u2606_o_placeOpt_3}),
    .c({_al_u2606_o_placeOpt_3,\t/a/reg_writedat [27]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aludat [27],open_n16693}),
    .e({\t/a/ID_read_dat2 [27],_al_u2610_o_placeOpt_3}),
    .mi({open_n16695,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [27],_al_u2631_o}),
    .q({open_n16710,\t/a/regfile/regfile$3$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2634 (
    .a({\t/a/aludat [27],\t/a/aludat [27]}),
    .b({_al_u2633_o,_al_u2633_o}),
    .c({_al_u2614_o_placeOpt_2,_al_u2614_o_placeOpt_2}),
    .d({_al_u2616_o_placeOpt_2,_al_u2616_o_placeOpt_2}),
    .mi({open_n16723,\t/a/ID_read_dat1 [27]}),
    .fx({open_n16728,\t/a/ID_jump_regdat1 [27]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(A*(C*~(1)*~(D)+C*1*~(D)+~(C)*1*D+C*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1110111011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2638 (
    .a({_al_u2614_o_placeOpt_2,\t/a/aludat [26]}),
    .b({_al_u2637_o,_al_u2637_o}),
    .c({\t/a/aludat [26],_al_u2614_o_placeOpt_2}),
    .d({_al_u2616_o_placeOpt_2,_al_u2616_o_placeOpt_2}),
    .mi({open_n16743,\t/a/ID_read_dat1 [26]}),
    .fx({open_n16748,\t/a/ID_jump_regdat1 [26]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2640 (
    .a({\t/a/aludat [25],\t/a/aludat [25]}),
    .b({_al_u2639_o,_al_u2639_o}),
    .c({_al_u2606_o,_al_u2606_o}),
    .d({_al_u2610_o,_al_u2610_o}),
    .mi({open_n16763,\t/a/ID_read_dat2 [25]}),
    .fx({open_n16768,\t/a/ID_jump_regdat2 [25]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~C*~A*~D+~B*~C*A*~D+~B*~C*~A*D+B*~C*~A*D+B*C*~A*D+~B*~C*A*D+B*~C*A*D+B*C*A*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("B*~C*~A*D+B*C*~A*D+B*~C*A*D+B*C*A*D"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b1110110011001100),
    .INIT_LUTG0(16'b1100110000000000),
    .INIT_LUTG1(16'b1111110011011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2642|t/a/id_ex/reg8_b25  (
    .a({_al_u2616_o_placeOpt_1,open_n16771}),
    .b({_al_u2641_o,_al_u333_o}),
    .c({_al_u2614_o_placeOpt_2,_al_u637_o}),
    .clk(clock_pad),
    .d({\t/a/ID_read_dat1 [25],\t/a/reg_writedat [25]}),
    .e({\t/a/aludat [25],_al_u647_o}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [25],\t/a/ID_read_dat1 [25]}),
    .q({open_n16790,\t/a/EX_regdat1 [25]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*~C*D+~B*A*~C*D+~B*~A*C*D+~B*A*C*D"),
    //.LUTF1("~(~A*~(C*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)))"),
    //.LUTG0("~B*~A*C*~D+~B*A*C*~D+~B*~A*C*D+~B*A*C*D"),
    //.LUTG1("~(~A*~(C*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100000000),
    .INIT_LUTF1(16'b1010101011101010),
    .INIT_LUTG0(16'b0011000000110000),
    .INIT_LUTG1(16'b1111101011101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2644|t/a/regfile/reg0_b120  (
    .a({_al_u2643_o,open_n16791}),
    .b({\t/a/aludat [24],_al_u2606_o_placeOpt_3}),
    .c({_al_u2606_o_placeOpt_3,\t/a/MEM_aludat [24]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o_placeOpt_3,\t/a/reg_writedat [24]}),
    .e({\t/a/ID_read_dat2 [24],_al_u2610_o_placeOpt_3}),
    .mi({open_n16793,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [24],_al_u2643_o}),
    .q({open_n16808,\t/a/regfile/regfile$3$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100000101),
    .INIT_LUTF1(16'b1110110011101100),
    .INIT_LUTG0(16'b1010101000000000),
    .INIT_LUTG1(16'b1111110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2646|t/a/id_ex/reg8_b24  (
    .a({\t/a/aludat [24],_al_u333_o}),
    .b({_al_u2645_o,open_n16809}),
    .c({_al_u2614_o_placeOpt_2,_al_u668_o}),
    .clk(clock_pad),
    .d({\t/a/ID_read_dat1 [24],\t/a/reg_writedat [24]}),
    .e({_al_u2616_o_placeOpt_2,_al_u658_o}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [24],\t/a/ID_read_dat1 [24]}),
    .q({open_n16828,\t/a/EX_regdat1 [24]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*B*A*~D+C*B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTF1("~(~A*~(C*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)))"),
    //.LUTG0("0"),
    //.LUTG1("~(~A*~(C*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101110001000),
    .INIT_LUTF1(16'b1010101011101010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111101011101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2648|t/a/regfile/reg0_b119  (
    .a({_al_u2647_o,\t/a/MEM_aludat [23]}),
    .b({\t/a/aludat [23],_al_u2610_o_placeOpt_3}),
    .c({_al_u2606_o_placeOpt_3,open_n16829}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o_placeOpt_3,\t/a/reg_writedat [23]}),
    .e({\t/a/ID_read_dat2 [23],_al_u2606_o_placeOpt_3}),
    .mi({open_n16831,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [23],_al_u2647_o}),
    .q({open_n16846,\t/a/regfile/regfile$3$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2652|_al_u2654  (
    .a({\t/a/aludat [22],\t/a/aludat [22]}),
    .b({_al_u2651_o,_al_u2653_o}),
    .c({_al_u2606_o_placeOpt_3,_al_u2614_o_placeOpt_2}),
    .d({_al_u2610_o_placeOpt_3,_al_u2616_o_placeOpt_2}),
    .e({\t/a/ID_read_dat2 [22],\t/a/ID_read_dat1 [22]}),
    .f({\t/a/ID_jump_regdat2 [22],\t/a/ID_jump_regdat1 [22]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2656 (
    .a({\t/a/aludat [21],\t/a/aludat [21]}),
    .b({_al_u2655_o,_al_u2655_o}),
    .c({_al_u2606_o_placeOpt_3,_al_u2606_o_placeOpt_3}),
    .d({_al_u2610_o_placeOpt_3,_al_u2610_o_placeOpt_3}),
    .mi({open_n16881,\t/a/ID_read_dat2 [21]}),
    .fx({open_n16886,\t/a/ID_jump_regdat2 [21]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~A*~C*~B+~D*A*~C*~B+~D*~A*~C*B+D*~A*~C*B+~D*A*~C*B+D*A*~C*B+D*~A*C*B+D*A*C*B"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("D*~A*~C*B+D*A*~C*B+D*~A*C*B+D*A*C*B"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100110000001111),
    .INIT_LUTF1(16'b1100110011001100),
    .INIT_LUTG0(16'b1100110000000000),
    .INIT_LUTG1(16'b1110111011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2658|t/a/id_ex/reg8_b21  (
    .a({\t/a/ID_read_dat1 [21],open_n16889}),
    .b({_al_u2657_o,\t/a/reg_writedat [21]}),
    .c({\t/a/aludat [21],_al_u731_o}),
    .clk(clock_pad),
    .d({_al_u2616_o_placeOpt_2,_al_u333_o}),
    .e({_al_u2614_o_placeOpt_2,_al_u721_o}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [21],\t/a/ID_read_dat1 [21]}),
    .q({open_n16908,\t/a/EX_regdat1 [21]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*D+~A*C*~B*D+~A*~C*B*D+~A*C*B*D"),
    //.LUTF1("~(~A*~(C*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)))"),
    //.LUTG0("~A*~C*B*~D+~A*C*B*~D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG1("~(~A*~(C*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010100000000),
    .INIT_LUTF1(16'b1010101011101010),
    .INIT_LUTG0(16'b0100010001000100),
    .INIT_LUTG1(16'b1111101011101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2660|t/a/regfile/reg0_b116  (
    .a({_al_u2659_o,_al_u2606_o_placeOpt_1}),
    .b({\t/a/aludat [20],\t/a/MEM_aludat [20]}),
    .c({_al_u2606_o_placeOpt_1,open_n16909}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o_placeOpt_1,\t/a/reg_writedat [20]}),
    .e({\t/a/ID_read_dat2 [20],_al_u2610_o_placeOpt_1}),
    .mi({open_n16911,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [20],_al_u2659_o}),
    .q({open_n16926,\t/a/regfile/regfile$3$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000011),
    .INIT_LUTF1(16'b1110110011101100),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1111110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2662|t/a/id_ex/reg8_b20  (
    .a({\t/a/aludat [20],open_n16927}),
    .b({_al_u2661_o,_al_u742_o}),
    .c({_al_u2614_o_placeOpt_2,_al_u752_o}),
    .clk(clock_pad),
    .d({\t/a/ID_read_dat1 [20],\t/a/reg_writedat [20]}),
    .e({_al_u2616_o_placeOpt_2,_al_u333_o}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [20],\t/a/ID_read_dat1 [20]}),
    .q({open_n16946,\t/a/EX_regdat1 [20]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~(~D*~(C*(B*~(0)*~(A)+B*0*~(A)+~(B)*0*A+B*0*A)))"),
    //.LUTG0("0"),
    //.LUTG1("~(~D*~(C*(B*~(1)*~(A)+B*1*~(A)+~(B)*1*A+B*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b1111111101000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111111111100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2664|t/a/regfile/reg0_b115  (
    .a({_al_u2610_o,open_n16947}),
    .b({\t/a/aludat [19],_al_u2610_o}),
    .c({_al_u2606_o,\t/a/MEM_aludat [19]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2663_o,\t/a/reg_writedat [19]}),
    .e({\t/a/ID_read_dat2 [19],_al_u2606_o}),
    .mi({open_n16949,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [19],_al_u2663_o}),
    .q({open_n16964,\t/a/regfile/regfile$3$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2666 (
    .a({\t/a/aludat [19],\t/a/aludat [19]}),
    .b({_al_u2665_o,_al_u2665_o}),
    .c({_al_u2614_o_placeOpt_2,_al_u2614_o_placeOpt_2}),
    .d({_al_u2616_o_placeOpt_2,_al_u2616_o_placeOpt_2}),
    .mi({open_n16977,\t/a/ID_read_dat1 [19]}),
    .fx({open_n16982,\t/a/ID_jump_regdat1 [19]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*~C*~A+~B*D*~C*~A+~B*~D*~C*A+B*~D*~C*A+~B*D*~C*A+B*D*~C*A+B*~D*C*A+B*D*C*A"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("B*~D*~C*A+B*D*~C*A+B*~D*C*A+B*D*C*A"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000101110001011),
    .INIT_LUTF1(16'b1110110011001100),
    .INIT_LUTG0(16'b1000100010001000),
    .INIT_LUTG1(16'b1110110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2670|t/a/id_ex/reg8_b18  (
    .a({\t/a/ID_read_dat1 [18],\t/a/reg_writedat [18]}),
    .b({_al_u2669_o,_al_u333_o}),
    .c({_al_u2614_o_placeOpt_2,_al_u815_o}),
    .clk(clock_pad),
    .d({_al_u2616_o_placeOpt_2,open_n16986}),
    .e({\t/a/aludat [18],_al_u805_o}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [18],\t/a/ID_read_dat1 [18]}),
    .q({open_n17004,\t/a/EX_regdat1 [18]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~D*~C+~A*~B*D*~C+~A*~B*~D*C+A*~B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+A*B*D*C"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("A*~B*~D*C+A*B*~D*C+A*~B*D*C+A*B*D*C"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000110110001),
    .INIT_LUTF1(16'b1110101011101010),
    .INIT_LUTG0(16'b1010000010100000),
    .INIT_LUTG1(16'b1111101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2674|t/a/id_ex/reg8_b17  (
    .a({_al_u2673_o,_al_u333_o}),
    .b({\t/a/aludat [17],_al_u826_o}),
    .c({_al_u2614_o_placeOpt_2,\t/a/reg_writedat [17]}),
    .clk(clock_pad),
    .d({\t/a/ID_read_dat1 [17],open_n17006}),
    .e({_al_u2616_o_placeOpt_2,_al_u836_o}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [17],\t/a/ID_read_dat1 [17]}),
    .q({open_n17024,\t/a/EX_regdat1 [17]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2676 (
    .a({\t/a/aludat [16],\t/a/aludat [16]}),
    .b({_al_u2675_o,_al_u2675_o}),
    .c({_al_u2606_o_placeOpt_3,_al_u2606_o_placeOpt_3}),
    .d({_al_u2610_o_placeOpt_3,_al_u2610_o_placeOpt_3}),
    .mi({open_n17037,\t/a/ID_read_dat2 [16]}),
    .fx({open_n17042,\t/a/ID_jump_regdat2 [16]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTF1("~(~D*~(A*(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("0"),
    //.LUTG1("~(~D*~(A*(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110001011100010),
    .INIT_LUTF1(16'b1111111100100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111111110101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2678|t/a/regfile/reg0_b1008  (
    .a({_al_u2614_o_placeOpt_2,\t/a/reg_writedat [16]}),
    .b({_al_u2616_o_placeOpt_1,_al_u2616_o_placeOpt_1}),
    .c({\t/a/aludat [16],\t/a/MEM_aludat [16]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2677_o,open_n17045}),
    .e({\t/a/ID_read_dat1 [16],_al_u2614_o_placeOpt_2}),
    .mi({open_n17047,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [16],_al_u2677_o}),
    .q({open_n17062,\t/a/regfile/regfile$31$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~D*~C+A*B*~D*~C+~A*B*D*~C+A*B*D*~C+~A*B*~D*C+~A*B*D*C"),
    //.LUTF1("A*C*~B*~D+A*C*B*~D+A*C*~B*D+A*C*B*D"),
    //.LUTG0("~A*B*~D*~C+A*B*~D*~C+~A*B*D*~C+A*B*D*~C"),
    //.LUTG1("~A*C*~B*~D+A*C*~B*~D+~A*C*B*~D+A*C*B*~D+~A*C*~B*D+A*C*~B*D+~A*C*B*D+A*C*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100110001001100),
    .INIT_LUTF1(16'b1010000010100000),
    .INIT_LUTG0(16'b0000110000001100),
    .INIT_LUTG1(16'b1111000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2679|t/a/ex_mem/reg4_b15  (
    .a({_al_u2427_o,_al_u2427_o}),
    .b({open_n17063,_al_u2435_o}),
    .c({_al_u2128_o,_al_u2128_o}),
    .clk(clock_pad),
    .e({_al_u2436_o,_al_u2436_o}),
    .sr(rst_pad),
    .f({_al_u2679_o,open_n17081}),
    .q({open_n17085,\t/a/MEM_aludat [15]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~A*C))"),
    //.LUT1("(D*~(~C*A))"),
    .INIT_LUT0(16'b1010111100000000),
    .INIT_LUT1(16'b1111010100000000),
    .MODE("LOGIC"))
    \_al_u2680|_al_u2748  (
    .a({_al_u2610_o,\t/a/ID_read_dat2 [3]}),
    .c({\t/a/ID_read_dat2 [15],_al_u2610_o}),
    .d({_al_u2606_o,_al_u2606_o}),
    .f({_al_u2680_o,_al_u2748_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(B*~A))))"),
    .INIT_LUT0(16'b1111111101000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2682 (
    .a({_al_u2679_o,_al_u2679_o}),
    .b({_al_u2435_o,_al_u2435_o}),
    .c({_al_u2680_o,_al_u2680_o}),
    .d({_al_u2681_o,_al_u2681_o}),
    .mi({open_n17120,_al_u2610_o_placeOpt_3}),
    .fx({open_n17125,\t/a/ID_jump_regdat2 [15]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~D*B+A*~C*~D*B+~A*~C*D*B+A*~C*D*B"),
    //.LUTF1("~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTG0("~A*~C*~D*B+A*~C*~D*B+~A*C*~D*B+A*C*~D*B+~A*~C*D*B+A*~C*D*B+~A*C*D*B+A*C*D*B"),
    //.LUTG1("~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    .INIT_LUTF0(16'b0000110000001100),
    .INIT_LUTF1(16'b1100110011001100),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b1100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2683|_al_u2713  (
    .b({_al_u2614_o_placeOpt_2,_al_u2614_o_placeOpt_2}),
    .c({\t/a/ID_read_dat1 [15],_al_u2616_o_placeOpt_1}),
    .e({_al_u2616_o_placeOpt_1,\t/a/ID_read_dat1 [10]}),
    .f({_al_u2683_o,_al_u2713_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*~C*A+~B*D*~C*A+~B*~D*C*A+~B*D*C*A"),
    //.LUTF1("~(~A*~(B*~(~0*~(C*~D))))"),
    //.LUTG0("~B*~D*C*~A+~B*D*C*~A+~B*~D*C*A+~B*D*C*A"),
    //.LUTG1("~(~A*~(B*~(~1*~(C*~D))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000100010),
    .INIT_LUTF1(16'b1010101011101010),
    .INIT_LUTG0(16'b0011000000110000),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2685|t/a/regfile/reg0_b1007  (
    .a({_al_u2684_o,\t/a/reg_writedat [15]}),
    .b({_al_u2683_o,_al_u2614_o_placeOpt_2}),
    .c({_al_u2435_o,\t/a/MEM_aludat [15]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2679_o,open_n17154}),
    .e({_al_u2616_o_placeOpt_2,_al_u2616_o_placeOpt_2}),
    .mi({open_n17156,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [15],_al_u2684_o}),
    .q({open_n17171,\t/a/regfile/regfile$31$ [15]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~(~0*A))"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*A*C*~D+B*A*C*~D"),
    //.LUTG0("(D*~C*~B*~(~1*A))"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0000000010101111),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2688|_al_u2687  (
    .a({\t/a/alu/n6 [14],\t/a/alu/n5 [14]}),
    .b({open_n17172,_al_u2686_o}),
    .c({_al_u2126_o,\t/a/EX_operation [2]}),
    .d({_al_u2687_o,_al_u2128_o}),
    .e({_al_u2439_o,\t/a/EX_operation$0$_lutinv_placeOpt_5 }),
    .f({_al_u2688_o,_al_u2687_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~A*C))"),
    //.LUT1("(D*~(~A*C))"),
    .INIT_LUT0(16'b1010111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"))
    \_al_u2690|_al_u2729  (
    .a({\t/a/ID_read_dat2 [14],\t/a/ID_read_dat2 [6]}),
    .c({_al_u2610_o,_al_u2610_o}),
    .d({_al_u2606_o,_al_u2606_o}),
    .f({_al_u2690_o,_al_u2729_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(~0*~(~B*A))))"),
    //.LUTF1("~(~C*~(D*~(~0*~(~B*A))))"),
    //.LUTG0("~(~D*~(C*~(~1*~(~B*A))))"),
    //.LUTG1("~(~C*~(D*~(~1*~(~B*A))))"),
    .INIT_LUTF0(16'b1111111100100000),
    .INIT_LUTF1(16'b1111001011110000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2691|_al_u2694  (
    .a({_al_u2688_o,_al_u2688_o}),
    .b({_al_u2446_o,_al_u2446_o}),
    .c({_al_u2689_o,_al_u2692_o}),
    .d({_al_u2690_o,_al_u2693_o}),
    .e({_al_u2610_o_placeOpt_1,_al_u2616_o_placeOpt_2}),
    .f({\t/a/ID_jump_regdat2 [14],\t/a/ID_jump_regdat1 [14]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2696 (
    .a({_al_u2610_o_placeOpt_3,\t/a/aludat [13]}),
    .b({_al_u2695_o,_al_u2695_o}),
    .c({_al_u2606_o_placeOpt_3,_al_u2606_o_placeOpt_3}),
    .d({\t/a/aludat [13],_al_u2610_o_placeOpt_3}),
    .mi({open_n17251,\t/a/ID_read_dat2 [13]}),
    .fx({open_n17256,\t/a/ID_jump_regdat2 [13]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(A*(C*~(1)*~(D)+C*1*~(D)+~(C)*1*D+C*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1110111011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2698 (
    .a({_al_u2614_o_placeOpt_2,\t/a/aludat [13]}),
    .b({_al_u2697_o,_al_u2697_o}),
    .c({\t/a/aludat [13],_al_u2614_o_placeOpt_2}),
    .d({_al_u2616_o_placeOpt_2,_al_u2616_o_placeOpt_2}),
    .mi({open_n17271,\t/a/ID_read_dat1 [13]}),
    .fx({open_n17276,\t/a/ID_jump_regdat1 [13]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*A*~C+D*B*A*~C+~D*~B*~A*C+D*~B*~A*C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTF1("~(~D*~(C*(B*~(0)*~(A)+B*0*~(A)+~(B)*0*A+B*0*A)))"),
    //.LUTG0("0"),
    //.LUTG1("~(~D*~(C*(B*~(1)*~(A)+B*1*~(A)+~(B)*1*A+B*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011100010111000),
    .INIT_LUTF1(16'b1111111101000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111111111100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2702|t/a/regfile/reg0_b1004  (
    .a({_al_u2616_o_placeOpt_2,\t/a/MEM_aludat [12]}),
    .b({\t/a/aludat [12],_al_u2616_o_placeOpt_2}),
    .c({_al_u2614_o_placeOpt_2,\t/a/reg_writedat [12]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2701_o,open_n17279}),
    .e({\t/a/ID_read_dat1 [12],_al_u2614_o_placeOpt_2}),
    .mi({open_n17281,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [12],_al_u2701_o}),
    .q({open_n17296,\t/a/regfile/regfile$31$ [12]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*~C*A+~B*D*~C*A+~B*~D*C*A+~B*D*C*A"),
    //.LUTF1("~(~D*~(C*(B*~(0)*~(A)+B*0*~(A)+~(B)*0*A+B*0*A)))"),
    //.LUTG0("~B*~D*C*~A+~B*D*C*~A+~B*~D*C*A+~B*D*C*A"),
    //.LUTG1("~(~D*~(C*(B*~(1)*~(A)+B*1*~(A)+~(B)*1*A+B*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000100010),
    .INIT_LUTF1(16'b1111111101000000),
    .INIT_LUTG0(16'b0011000000110000),
    .INIT_LUTG1(16'b1111111111100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2706|t/a/regfile/reg0_b1003  (
    .a({_al_u2616_o_placeOpt_2,\t/a/reg_writedat [11]}),
    .b({\t/a/aludat [11],_al_u2614_o_placeOpt_2}),
    .c({_al_u2614_o_placeOpt_2,\t/a/MEM_aludat [11]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2705_o,open_n17297}),
    .e({\t/a/ID_read_dat1 [11],_al_u2616_o_placeOpt_2}),
    .mi({open_n17299,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [11],_al_u2705_o}),
    .q({open_n17314,\t/a/regfile/regfile$31$ [11]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2708 (
    .a({\t/a/alu/n5 [10],\t/a/alu/n5 [10]}),
    .b({_al_u2707_o,_al_u2707_o}),
    .c({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n17327,\t/a/EX_operation$0$_lutinv_placeOpt_2 }),
    .fx({open_n17332,_al_u2708_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(~0*~(~B*A))))"),
    //.LUTF1("~(~D*~(C*~(~0*~(~B*A))))"),
    //.LUTG0("~(~D*~(C*~(~1*~(~B*A))))"),
    //.LUTG1("~(~D*~(C*~(~1*~(~B*A))))"),
    .INIT_LUTF0(16'b1111111100100000),
    .INIT_LUTF1(16'b1111111100100000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2712|_al_u2715  (
    .a({_al_u2709_o,_al_u2709_o}),
    .b({_al_u2486_o,_al_u2486_o}),
    .c({_al_u2710_o,_al_u2713_o}),
    .d({_al_u2711_o,_al_u2714_o}),
    .e({_al_u2610_o_placeOpt_1,_al_u2616_o_placeOpt_2}),
    .f({\t/a/ID_jump_regdat2 [10],\t/a/ID_jump_regdat1 [10]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(A*(C*~(1)*~(D)+C*1*~(D)+~(C)*1*D+C*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1110111011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2717 (
    .a({_al_u2606_o,\t/a/aludat [9]}),
    .b({_al_u2716_o,_al_u2716_o}),
    .c({\t/a/aludat [9],_al_u2606_o}),
    .d({_al_u2610_o,_al_u2610_o}),
    .mi({open_n17369,\t/a/ID_read_dat2 [9]}),
    .fx({open_n17374,\t/a/ID_jump_regdat2 [9]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2719|_al_u1065  (
    .a({\t/a/aludat [9],\t/a/ID_rs2$0$_placeOpt_19 }),
    .b({_al_u2718_o,\t/a/ID_rs2$1$_placeOpt_19 }),
    .c({_al_u2614_o_placeOpt_3,\t/a/ID_rs2$2$_placeOpt_6 }),
    .d({_al_u2616_o_placeOpt_1,\t/a/regfile/regfile$31$ [9]}),
    .e({\t/a/ID_read_dat1 [9],\t/a/regfile/regfile$30$ [9]}),
    .f({\t/a/ID_jump_regdat1 [9],_al_u1065_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~D*~A*C+~B*D*~A*C+~B*~D*A*C+~B*D*A*C"),
    //.LUTF1("~(~D*~(C*(A*~(0)*~(B)+A*0*~(B)+~(A)*0*B+A*0*B)))"),
    //.LUTG0("~B*~D*A*~C+~B*D*A*~C+~B*~D*A*C+~B*D*A*C"),
    //.LUTG1("~(~D*~(C*(A*~(1)*~(B)+A*1*~(B)+~(A)*1*B+A*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000000110000),
    .INIT_LUTF1(16'b1111111100100000),
    .INIT_LUTG0(16'b0010001000100010),
    .INIT_LUTG1(16'b1111111111100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2721|t/a/regfile/reg0_b136  (
    .a({\t/a/aludat [8],\t/a/MEM_aludat [8]}),
    .b({_al_u2610_o_placeOpt_1,_al_u2606_o_placeOpt_1}),
    .c({_al_u2606_o_placeOpt_1,\t/a/reg_writedat [8]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2720_o,open_n17399}),
    .e({\t/a/ID_read_dat2 [8],_al_u2610_o_placeOpt_1}),
    .mi({open_n17401,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [8],_al_u2720_o}),
    .q({open_n17416,\t/a/regfile/regfile$4$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000011),
    .INIT_LUTF1(16'b1110110011101100),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1111110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2723|t/a/id_ex/reg8_b8  (
    .a({\t/a/aludat [8],open_n17417}),
    .b({_al_u2722_o,_al_u364_o}),
    .c({_al_u2614_o_placeOpt_2,_al_u374_o}),
    .clk(clock_pad),
    .d({\t/a/ID_read_dat1 [8],\t/a/reg_writedat [8]}),
    .e({_al_u2616_o_placeOpt_2,_al_u333_o}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [8],\t/a/ID_read_dat1 [8]}),
    .q({open_n17436,\t/a/EX_regdat1 [8]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*B*A*~C+D*B*A*~C+~D*~B*~A*C+D*~B*~A*C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTF1("~(~A*~(C*(B*~(0)*~(D)+B*0*~(D)+~(B)*0*D+B*0*D)))"),
    //.LUTG0("0"),
    //.LUTG1("~(~A*~(C*(B*~(1)*~(D)+B*1*~(D)+~(B)*1*D+B*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011100010111000),
    .INIT_LUTF1(16'b1010101011101010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111101011101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2725|t/a/regfile/reg0_b135  (
    .a({_al_u2724_o,\t/a/MEM_aludat [7]}),
    .b({\t/a/aludat [7],_al_u2610_o_placeOpt_1}),
    .c({_al_u2606_o_placeOpt_1,\t/a/reg_writedat [7]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o_placeOpt_1,open_n17437}),
    .e({\t/a/ID_read_dat2 [7],_al_u2606_o_placeOpt_1}),
    .mi({open_n17439,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [7],_al_u2724_o}),
    .q({open_n17454,\t/a/regfile/regfile$4$ [7]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+~A*~C*B*~D+~A*~C*~B*D+A*~C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+A*C*B*D"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("A*~C*~B*D+A*C*~B*D+A*~C*B*D+A*C*B*D"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100000101),
    .INIT_LUTF1(16'b1110110011101100),
    .INIT_LUTG0(16'b1010101000000000),
    .INIT_LUTG1(16'b1111110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2727|t/a/id_ex/reg8_b7  (
    .a({\t/a/aludat [7],_al_u333_o}),
    .b({_al_u2726_o,open_n17455}),
    .c({_al_u2614_o_placeOpt_1,_al_u385_o}),
    .clk(clock_pad),
    .d({\t/a/ID_read_dat1 [7],\t/a/reg_writedat [7]}),
    .e({_al_u2616_o_placeOpt_2,_al_u395_o}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [7],\t/a/ID_read_dat1 [7]}),
    .q({open_n17474,\t/a/EX_regdat1 [7]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUTF1("~(~B*~(C*~(~0*~(D*~A))))"),
    //.LUTG0("~(~D*~(C*~(~1*~(B*~A))))"),
    //.LUTG1("~(~B*~(C*~(~1*~(D*~A))))"),
    .INIT_LUTF0(16'b1111111101000000),
    .INIT_LUTF1(16'b1101110011001100),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2731|_al_u2734  (
    .a({_al_u2728_o,_al_u2728_o}),
    .b({_al_u2730_o,_al_u2525_o}),
    .c({_al_u2729_o,_al_u2732_o}),
    .d({_al_u2525_o,_al_u2733_o}),
    .e({_al_u2610_o_placeOpt_1,_al_u2616_o_placeOpt_2}),
    .f({\t/a/ID_jump_regdat2 [6],\t/a/ID_jump_regdat1 [6]}));
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(C*~(~A*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1011000010110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2732|t/a/id_ex/reg8_b6  (
    .a({\t/a/ID_read_dat1 [6],_al_u333_o}),
    .b({_al_u2616_o_placeOpt_1,_al_u406_o}),
    .c({_al_u2614_o_placeOpt_2,_al_u416_o}),
    .clk(clock_pad),
    .d({open_n17498,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u2732_o,\t/a/ID_read_dat1 [6]}),
    .q({open_n17514,\t/a/EX_regdat1 [6]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(~(A)*~(B)*~(D)+~(A)*~(B)*D+A*~(B)*D+~(A)*B*D))"),
    //.LUT1("(B*~(~D*~(~C*~A)))"),
    .INIT_LUT0(16'b0111000000010000),
    .INIT_LUT1(16'b1100110000000100),
    .MODE("LOGIC"))
    \_al_u2735|_al_u2536  (
    .a({\t/a/alu/mux0_b5/B1_0 ,\t/a/EX_A [5]}),
    .b({_al_u2128_o,\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o }),
    .c(\t/a/EX_operation [2:1]),
    .d({_al_u2536_o,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .f({_al_u2735_o,_al_u2536_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(A*~(~0*~(B*~C))))"),
    //.LUTF1("(A*~(~C*B))"),
    //.LUTG0("~(~D*~(A*~(~1*~(B*~C))))"),
    //.LUTG1("(A*~(~C*B))"),
    .INIT_LUTF0(16'b1111111100001000),
    .INIT_LUTF1(16'b1010001010100010),
    .INIT_LUTG0(16'b1111111110101010),
    .INIT_LUTG1(16'b1010001010100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2736|_al_u2738  (
    .a({_al_u2606_o_placeOpt_1,_al_u2736_o}),
    .b({_al_u2610_o_placeOpt_1,_al_u2535_o}),
    .c({\t/a/ID_read_dat2 [5],_al_u2735_o}),
    .d({open_n17537,_al_u2737_o}),
    .e({open_n17538,_al_u2610_o_placeOpt_1}),
    .f({_al_u2736_o,\t/a/ID_jump_regdat2 [5]}));
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(D*~(~A*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1011101100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2739|t/a/id_ex/reg8_b5  (
    .a({\t/a/ID_read_dat1 [5],_al_u333_o}),
    .b({_al_u2616_o_placeOpt_1,_al_u427_o}),
    .c({open_n17559,_al_u437_o}),
    .clk(clock_pad),
    .d({_al_u2614_o_placeOpt_3,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u2739_o,\t/a/ID_read_dat1 [5]}),
    .q({open_n17576,\t/a/EX_regdat1 [5]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(B*~A))))"),
    .INIT_LUT0(16'b1111111101000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2741 (
    .a({_al_u2735_o,_al_u2735_o}),
    .b({_al_u2535_o,_al_u2535_o}),
    .c({_al_u2739_o,_al_u2739_o}),
    .d({_al_u2740_o,_al_u2740_o}),
    .mi({open_n17589,_al_u2616_o_placeOpt_2}),
    .fx({open_n17594,\t/a/ID_jump_regdat1 [5]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2743 (
    .a({\t/a/aludat [4],\t/a/aludat [4]}),
    .b({_al_u2742_o,_al_u2742_o}),
    .c({_al_u2606_o_placeOpt_1,_al_u2606_o_placeOpt_1}),
    .d({_al_u2610_o_placeOpt_1,_al_u2610_o_placeOpt_1}),
    .mi({open_n17609,\t/a/ID_read_dat2 [4]}),
    .fx({open_n17614,\t/a/ID_jump_regdat2 [4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~C*~A*~D+~B*~C*A*~D+~B*~C*~A*D+B*~C*~A*D+B*C*~A*D+~B*~C*A*D+B*~C*A*D+B*C*A*D"),
    //.LUTF1("~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTG0("B*~C*~A*D+B*C*~A*D+B*~C*A*D+B*C*A*D"),
    //.LUTG1("A*~D*~C*B+A*D*~C*B+A*~D*C*B+A*D*C*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111100000011),
    .INIT_LUTF1(16'b1100110011001100),
    .INIT_LUTG0(16'b1100110000000000),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2744|t/a/id_ex/reg8_b4  (
    .a({\t/a/ID_read_dat1 [4],open_n17617}),
    .b({_al_u2614_o,_al_u333_o}),
    .c({open_n17618,_al_u448_o}),
    .clk(clock_pad),
    .d({open_n17620,\t/a/reg_writedat [4]}),
    .e({_al_u2616_o,_al_u458_o}),
    .sr(rst_pad),
    .f({_al_u2744_o,\t/a/ID_read_dat1 [4]}),
    .q({open_n17638,\t/a/EX_regdat1 [4]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("~(~A*~((~B*~C))*~(D)+~A*(~B*~C)*~(D)+~(~A)*(~B*~C)*D+~A*(~B*~C)*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b1111110010101010),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2746|t/a/regfile/reg0_b132  (
    .a({_al_u2745_o,_al_u2614_o_placeOpt_1}),
    .b({\t/a/aludat [4],_al_u2616_o_placeOpt_2}),
    .c({_al_u2616_o_placeOpt_2,\t/a/MEM_aludat [4]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2744_o,\t/a/reg_writedat [4]}),
    .mi({open_n17649,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [4],_al_u2745_o}),
    .q({open_n17653,\t/a/regfile/regfile$4$ [4]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(~(A)*~(B)*~(D)+~(A)*~(B)*D+A*~(B)*D+~(A)*B*D))"),
    //.LUT1("(A*~(~D*~(~C*~B)))"),
    .INIT_LUT0(16'b0111000000010000),
    .INIT_LUT1(16'b1010101000000010),
    .MODE("LOGIC"))
    \_al_u2747|_al_u2556  (
    .a({_al_u2128_o,\t/a/EX_A [3]}),
    .b({\t/a/alu/mux0_b3/B1_0 ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_4 }),
    .c(\t/a/EX_operation [2:1]),
    .d({_al_u2556_o,\t/a/EX_operation$0$_lutinv_placeOpt_1 }),
    .f({_al_u2747_o,_al_u2556_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(B*~A))))"),
    .INIT_LUT0(16'b1111111101000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2750 (
    .a({_al_u2747_o,_al_u2747_o}),
    .b({_al_u2555_o,_al_u2555_o}),
    .c({_al_u2748_o,_al_u2748_o}),
    .d({_al_u2749_o,_al_u2749_o}),
    .mi({open_n17686,_al_u2610_o_placeOpt_3}),
    .fx({open_n17691,\t/a/ID_jump_regdat2 [3]}));
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(D*~(~A*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2751|t/a/id_ex/reg8_b3  (
    .a({\t/a/ID_read_dat1 [3],_al_u333_o}),
    .b({open_n17694,_al_u469_o}),
    .c({_al_u2616_o_placeOpt_3,_al_u479_o}),
    .clk(clock_pad),
    .d({_al_u2614_o,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u2751_o,\t/a/ID_read_dat1 [3]}),
    .q({open_n17711,\t/a/EX_regdat1 [3]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(B*~A))))"),
    .INIT_LUT0(16'b1111111101000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2753 (
    .a({_al_u2747_o,_al_u2747_o}),
    .b({_al_u2555_o,_al_u2555_o}),
    .c({_al_u2751_o,_al_u2751_o}),
    .d({_al_u2752_o,_al_u2752_o}),
    .mi({open_n17724,_al_u2616_o_placeOpt_2}),
    .fx({open_n17729,\t/a/ID_jump_regdat1 [3]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2755|_al_u2757  (
    .a({\t/a/aludat [2],\t/a/aludat [2]}),
    .b({_al_u2754_o,_al_u2756_o}),
    .c({_al_u2606_o_placeOpt_1,_al_u2614_o_placeOpt_1}),
    .d({_al_u2610_o_placeOpt_1,_al_u2616_o_placeOpt_2}),
    .e({\t/a/ID_read_dat2 [2],\t/a/ID_read_dat1 [2]}),
    .f({\t/a/ID_jump_regdat2 [2],\t/a/ID_jump_regdat1 [2]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2759|_al_u2761  (
    .a({\t/a/aludat [0],\t/a/aludat [0]}),
    .b({_al_u2758_o,_al_u2760_o}),
    .c({_al_u2606_o_placeOpt_1,_al_u2614_o_placeOpt_1}),
    .d({_al_u2610_o_placeOpt_1,_al_u2616_o_placeOpt_2}),
    .e({\t/a/ID_read_dat2 [0],\t/a/ID_read_dat1 [0]}),
    .f({\t/a/ID_jump_regdat2 [0],\t/a/ID_jump_regdat1 [0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*~A)"),
    //.LUT1("(~1*~D*~A*~B*~C)"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u276 (
    .a({\t/a/WB_rd [2],\t/a/WB_rd [0]}),
    .b({\t/a/WB_rd [1],\t/a/WB_rd [1]}),
    .c({\t/a/WB_rd [0],\t/a/WB_rd [2]}),
    .d({\t/a/WB_rd [3],\t/a/WB_rd [3]}),
    .mi({open_n17788,\t/a/WB_rd [4]}),
    .fx({open_n17793,\t/a/regfile/n46 [0]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~(~D*~(A*(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("~(~D*~(A*(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010100000000),
    .INIT_LUTF1(16'b1111111100100000),
    .INIT_LUTG0(16'b0101000001010000),
    .INIT_LUTG1(16'b1111111110101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2763|t/a/regfile/reg0_b129  (
    .a({_al_u2606_o_placeOpt_1,_al_u2606_o_placeOpt_1}),
    .b({_al_u2610_o_placeOpt_1,open_n17796}),
    .c({\t/a/aludat [1],\t/a/MEM_aludat [1]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2762_o,\t/a/reg_writedat [1]}),
    .e({\t/a/ID_read_dat2 [1],_al_u2610_o_placeOpt_1}),
    .mi({open_n17798,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [1],_al_u2762_o}),
    .q({open_n17813,\t/a/regfile/regfile$4$ [1]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2765 (
    .a({\t/a/aludat [1],\t/a/aludat [1]}),
    .b({_al_u2764_o,_al_u2764_o}),
    .c({_al_u2614_o_placeOpt_1,_al_u2614_o_placeOpt_1}),
    .d({_al_u2616_o_placeOpt_2,_al_u2616_o_placeOpt_2}),
    .mi({open_n17826,\t/a/ID_read_dat1 [1]}),
    .fx({open_n17831,\t/a/ID_jump_regdat1 [1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~A*~C*~B+D*A*~C*~B+~D*~A*C*~B+D*A*C*~B+~D*~A*~C*B+D*A*~C*B+~D*~A*C*B+D*A*C*B"),
    //.LUTF1("~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG0("~D*~A*C*~B+D*A*C*~B+~D*~A*C*B+D*A*C*B"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1010101001010101),
    .INIT_LUTF1(16'b1111000011110000),
    .INIT_LUTG0(16'b1010000001010000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2767|_al_u2770  (
    .a({open_n17834,\t/a/ID_jump_regdat1 [14]}),
    .c({\t/a/ID_jump_regdat2 [1],\t/a/ID_jump_regdat2 [1]}),
    .d({open_n17839,\t/a/ID_jump_regdat2 [14]}),
    .e({\t/a/ID_jump_regdat1 [1],\t/a/ID_jump_regdat1 [1]}),
    .f({_al_u2767_o,_al_u2770_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0@D)*~(C@B))"),
    //.LUT1("(~A*~(1@D)*~(C@B))"),
    .INIT_LUT0(16'b0000000001000001),
    .INIT_LUT1(16'b0100000100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2768 (
    .a({_al_u2767_o,_al_u2767_o}),
    .b({\t/a/ID_jump_regdat2 [13],\t/a/ID_jump_regdat2 [13]}),
    .c({\t/a/ID_jump_regdat1 [13],\t/a/ID_jump_regdat1 [13]}),
    .d({\t/a/ID_jump_regdat2 [4],\t/a/ID_jump_regdat2 [4]}),
    .mi({open_n17872,\t/a/ID_jump_regdat1 [4]}),
    .fx({open_n17877,_al_u2768_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("~A*~B*~C*~D+A*B*~C*~D+~A*~B*C*D+A*B*C*D"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("~A*~B*~C*~D+A*B*~C*~D+~A*~B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1001000000001001),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1001000000001001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2769|_al_u2668  (
    .a({\t/a/ID_jump_regdat2 [18],\t/a/aludat [18]}),
    .b({\t/a/ID_jump_regdat1 [18],_al_u2667_o}),
    .c({\t/a/ID_jump_regdat1 [5],_al_u2606_o_placeOpt_1}),
    .d({\t/a/ID_jump_regdat2 [5],_al_u2610_o_placeOpt_1}),
    .e({open_n17882,\t/a/ID_read_dat2 [18]}),
    .f({_al_u2769_o,\t/a/ID_jump_regdat2 [18]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~C)*~(B*~A))"),
    //.LUT1("(~(D@C)*~(B@A))"),
    .INIT_LUT0(16'b1011000010111011),
    .INIT_LUT1(16'b1001000000001001),
    .MODE("LOGIC"))
    \_al_u2772|_al_u2776  (
    .a({\t/a/ID_jump_regdat2 [22],\t/a/ID_jump_regdat2 [28]}),
    .b({\t/a/ID_jump_regdat1 [22],\t/a/ID_jump_regdat1 [28]}),
    .c({\t/a/ID_jump_regdat2 [21],\t/a/ID_jump_regdat2 [26]}),
    .d({\t/a/ID_jump_regdat1 [21],\t/a/ID_jump_regdat1 [26]}),
    .f({_al_u2772_o,_al_u2776_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("0"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("A*~C*~D*~B+A*C*~D*~B+A*~C*D*B+A*C*D*B"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000100000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2773|_al_u2771  (
    .a({_al_u2771_o,_al_u2768_o}),
    .b({\t/a/ID_jump_regdat1 [31],_al_u2769_o}),
    .c({open_n17923,_al_u2770_o}),
    .d({\t/a/ID_jump_regdat2 [31],\t/a/ID_jump_regdat2 [10]}),
    .e({_al_u2772_o,\t/a/ID_jump_regdat1 [10]}),
    .f({_al_u2773_o,_al_u2771_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("(~B*D)"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("(~B*D)"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b0011001100000000),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b0011001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2774|_al_u2636  (
    .a({open_n17946,\t/a/aludat [26]}),
    .b({\t/a/ID_jump_regdat1 [26],_al_u2635_o}),
    .c({open_n17947,_al_u2606_o_placeOpt_3}),
    .d({\t/a/ID_jump_regdat2 [26],_al_u2610_o_placeOpt_3}),
    .e({open_n17950,\t/a/ID_read_dat2 [26]}),
    .f({_al_u2774_o,\t/a/ID_jump_regdat2 [26]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@D)*~(~C*B))"),
    //.LUTF1("0"),
    //.LUTG0("(~A*~(1@D)*~(~C*B))"),
    //.LUTG1("B*A*~C*~D+B*A*C*D"),
    .INIT_LUTF0(16'b0000000001010001),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0101000100000000),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2777|_al_u2775  (
    .a({_al_u2775_o,_al_u2774_o}),
    .b({_al_u2773_o,\t/a/ID_jump_regdat2 [28]}),
    .c({\t/a/ID_jump_regdat2 [19],\t/a/ID_jump_regdat1 [28]}),
    .d({\t/a/ID_jump_regdat1 [19],\t/a/ID_jump_regdat2 [24]}),
    .e({_al_u2776_o,\t/a/ID_jump_regdat1 [24]}),
    .f({_al_u2777_o,_al_u2775_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("(~(C@D)*~(B@A))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("(~(C@D)*~(B@A))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1001000000001001),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1001000000001001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2778|_al_u2620  (
    .a({\t/a/ID_jump_regdat2 [30],\t/a/aludat [30]}),
    .b({\t/a/ID_jump_regdat1 [30],_al_u2619_o}),
    .c({\t/a/ID_jump_regdat1 [25],_al_u2606_o_placeOpt_3}),
    .d({\t/a/ID_jump_regdat2 [25],_al_u2610_o_placeOpt_3}),
    .e({open_n17995,\t/a/ID_read_dat2 [30]}),
    .f({_al_u2778_o,\t/a/ID_jump_regdat2 [30]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("A*~B*~C*~D+A*~B*C*D"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("A*B*~C*~D+A*B*C*D"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b0010000000000010),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2779|_al_u2624  (
    .a({_al_u2778_o,\t/a/aludat [29]}),
    .b({\t/a/ID_jump_regdat2 [29],_al_u2623_o}),
    .c({\t/a/ID_jump_regdat1 [27],_al_u2606_o_placeOpt_3}),
    .d({\t/a/ID_jump_regdat2 [27],_al_u2610_o_placeOpt_3}),
    .e({\t/a/ID_jump_regdat1 [29],\t/a/ID_read_dat2 [29]}),
    .f({_al_u2779_o,\t/a/ID_jump_regdat2 [29]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+A*~C*~B*~D+A*C*~B*~D+~A*~C*B*~D+A*~C*B*~D+A*C*B*~D"),
    //.LUTF1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~C*~B*D+A*~C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+A*C*B*D"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b0000000010101111),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b1010111100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2780|_al_u2782  (
    .a({open_n18038,\t/a/ID_jump_regdat2 [6]}),
    .c({open_n18041,\t/a/ID_jump_regdat1 [6]}),
    .d({\t/a/ID_jump_regdat2 [6],\t/a/ID_jump_regdat1 [2]}),
    .e({\t/a/ID_jump_regdat1 [6],\t/a/ID_jump_regdat2 [2]}),
    .f({_al_u2780_o,_al_u2782_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("~A*B*~C*~D+~A*B*C*D"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b0101000000000101),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b0100000000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2781|_al_u2672  (
    .a({_al_u2780_o,\t/a/aludat [17]}),
    .b({\t/a/ID_jump_regdat2 [20],_al_u2671_o}),
    .c({\t/a/ID_jump_regdat1 [17],_al_u2606_o_placeOpt_3}),
    .d({\t/a/ID_jump_regdat2 [17],_al_u2610_o_placeOpt_3}),
    .e({\t/a/ID_jump_regdat1 [20],\t/a/ID_read_dat2 [17]}),
    .f({_al_u2781_o,\t/a/ID_jump_regdat2 [17]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("0"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("~B*A*~C*~D+B*A*~C*~D+~B*A*C*D+B*A*C*D"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1010000000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2783|_al_u2650  (
    .a({_al_u2782_o,\t/a/aludat [23]}),
    .b({open_n18086,_al_u2649_o}),
    .c({\t/a/ID_jump_regdat1 [23],_al_u2614_o_placeOpt_2}),
    .d({\t/a/ID_jump_regdat2 [23],_al_u2616_o_placeOpt_2}),
    .e({_al_u2781_o,\t/a/ID_read_dat1 [23]}),
    .f({_al_u2783_o,\t/a/ID_jump_regdat1 [23]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("~A*~C*~B*~D+~A*C*~B*~D+~A*~C*B*D+~A*C*B*D"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("A*~C*~B*~D+A*C*~B*~D+A*~C*B*D+A*C*B*D"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b0100010000010001),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1000100000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2784|_al_u2700  (
    .a({\t/a/ID_jump_regdat2 [12],\t/a/aludat [12]}),
    .b({\t/a/ID_jump_regdat2 [8],_al_u2699_o}),
    .c({open_n18109,_al_u2606_o_placeOpt_3}),
    .d({\t/a/ID_jump_regdat1 [8],_al_u2610_o_placeOpt_3}),
    .e({\t/a/ID_jump_regdat1 [12],\t/a/ID_read_dat2 [12]}),
    .f({_al_u2784_o,\t/a/ID_jump_regdat2 [12]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(0@D)*~(C@B))"),
    //.LUT1("(A*~(1@B)*~(C@D))"),
    .INIT_LUT0(16'b0000000010000010),
    .INIT_LUT1(16'b1000000000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2787 (
    .a({_al_u2786_o,_al_u2786_o}),
    .b({\t/a/ID_jump_regdat2 [9],\t/a/ID_jump_regdat2 [0]}),
    .c({\t/a/ID_jump_regdat1 [0],\t/a/ID_jump_regdat1 [0]}),
    .d({\t/a/ID_jump_regdat2 [0],\t/a/ID_jump_regdat2 [9]}),
    .mi({open_n18144,\t/a/ID_jump_regdat1 [9]}),
    .fx({open_n18149,_al_u2787_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D@C)*~(~B*A))"),
    //.LUT1("(D*~C)"),
    .INIT_LUT0(16'b1101000000001101),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2788|_al_u2786  (
    .a({open_n18152,\t/a/ID_jump_regdat2 [15]}),
    .b({open_n18153,\t/a/ID_jump_regdat1 [15]}),
    .c({\t/a/ID_jump_regdat2 [15],\t/a/ID_jump_regdat2 [7]}),
    .d({\t/a/ID_jump_regdat1 [15],\t/a/ID_jump_regdat1 [7]}),
    .f({_al_u2788_o,_al_u2786_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("~A*~B*~C*~D+~A*~B*C*D"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("~A*B*~C*~D+~A*B*C*D"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b0001000000000001),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b0100000000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2789|_al_u2704  (
    .a({_al_u2788_o,\t/a/aludat [11]}),
    .b({\t/a/ID_jump_regdat2 [11],_al_u2703_o}),
    .c({\t/a/ID_jump_regdat2 [3],_al_u2606_o_placeOpt_3}),
    .d({\t/a/ID_jump_regdat1 [3],_al_u2610_o_placeOpt_3}),
    .e({\t/a/ID_jump_regdat1 [11],\t/a/ID_read_dat2 [11]}),
    .f({_al_u2789_o,\t/a/ID_jump_regdat2 [11]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0@D)*~(~C*B))"),
    //.LUTF1("(0*D*A*B*C)"),
    //.LUTG0("(A*~(1@D)*~(~C*B))"),
    //.LUTG1("(1*D*A*B*C)"),
    .INIT_LUTF0(16'b0000000010100010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010001000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2790|_al_u2785  (
    .a({_al_u2785_o,_al_u2784_o}),
    .b({_al_u2783_o,\t/a/ID_jump_regdat2 [20]}),
    .c({_al_u2779_o,\t/a/ID_jump_regdat1 [20]}),
    .d({_al_u2787_o,\t/a/ID_jump_regdat2 [16]}),
    .e({_al_u2789_o,\t/a/ID_jump_regdat1 [16]}),
    .f({_al_u2790_o,_al_u2785_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("~A*~C*~D*~B+A*~C*~D*~B+~A*C*~D*~B+A*C*~D*~B+~A*~C*D*~B+~A*C*D*~B"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("~A*~C*~D*~B+A*~C*~D*~B+~A*C*~D*~B+A*C*~D*~B"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0001000100110011),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2792|_al_u1756  (
    .a({_al_u2766_o,\t/a/condition/n5 [4]}),
    .b({\t/a/condition/sel1/B2 ,\t/a/condition/n0_lutinv }),
    .c({open_n18218,\t/a/condition/n1_lutinv }),
    .d({\t/a/condition/n1_lutinv ,\t/a/condition/sel1/B2 }),
    .e({_al_u2791_o,\t/a/ID_rd [4]}),
    .f({_al_u2792_o,\t/a/ID_jump_addr [4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+~A*B*C*D"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0101000011110000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0101010111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2794|_al_u1782  (
    .a({_al_u1958_o,\t/a/condition/n5 [1]}),
    .b({open_n18241,\t/a/condition/n0_lutinv }),
    .c({\t/a/ID_rd [1],\t/a/condition/n1_lutinv }),
    .d({\t/a/ID_rd [3],\t/a/condition/sel1/B2 }),
    .e({_al_u1965_o,\t/a/ID_rd [1]}),
    .f({_al_u2794_o,\t/a/ID_jump_addr [1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("~A*D*~C*~B+A*D*~C*~B+~A*D*C*~B+~A*D*~C*B+A*D*~C*B+~A*D*C*B"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+~A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+~A*D*C*B"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0101111100000000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0101111101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2795|_al_u1760  (
    .a({_al_u1962_o,\t/a/condition/n5 [3]}),
    .b({open_n18264,\t/a/condition/n0_lutinv }),
    .c({\t/a/ID_rd [0],\t/a/condition/n1_lutinv }),
    .d({_al_u1958_o,\t/a/condition/sel1/B2 }),
    .e({\t/a/ID_rd [3],\t/a/ID_rd [3]}),
    .f({_al_u2795_o,\t/a/ID_jump_addr [3]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(~C*B))"),
    //.LUT1("(~(B*D)*~(~A*~C))"),
    .INIT_LUT0(16'b1010111010101110),
    .INIT_LUT1(16'b0011001011111010),
    .MODE("LOGIC"))
    \_al_u2796|_al_u2091  (
    .a({\t/a/ID_rd [0],_al_u2078_o}),
    .b({\t/a/ID_rd [1],_al_u2080_o}),
    .c({_al_u1962_o,_al_u1962_o}),
    .d({_al_u1965_o,open_n18289}),
    .f({_al_u2796_o,\t/a/IF_skip_addr [20]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~B)"),
    //.LUTF1("0"),
    //.LUTG0("(A*~B)"),
    //.LUTG1("~B*C*A*D+B*C*A*D"),
    .INIT_LUTF0(16'b0010001000100010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0010001000100010),
    .INIT_LUTG1(16'b1010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2797|_al_u1742  (
    .a({_al_u2795_o,\t/a/ID_rs1$2$_placeOpt_10 }),
    .b({open_n18308,\t/a/EX_rd [2]}),
    .c({_al_u2794_o,open_n18309}),
    .d({_al_u2796_o,open_n18312}),
    .e({_al_u2793_o,open_n18313}),
    .f({\t/a/n4_lutinv ,_al_u1742_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("A*~C*~B*D+~A*C*~B*D+A*C*~B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111101000000000),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b1111101011111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2798|t/a/id_ex/reg5_b1  (
    .a({_al_u2113_o,open_n18334}),
    .b({open_n18335,\t/a/ID_rd [1]}),
    .c({\t/a/ID_rd [3],open_n18336}),
    .clk(clock_pad),
    .d({_al_u2117_o,open_n18338}),
    .e({\t/a/ID_rd [1],_al_u2117_o}),
    .mi({open_n18340,\t/a/ID_rd [1]}),
    .sr(rst_pad),
    .f({_al_u2798_o,_al_u2800_o}),
    .q({open_n18355,\t/a/EX_rd [1]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~A)"),
    //.LUT1("(D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b1010101000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2802|t/a/if_id/reg6_b3  (
    .a({\t/instruction$2$_neg_lutinv ,\t/a/if_id/n9 }),
    .clk(clock_pad),
    .d({\t/instruction$3$_neg_lutinv ,\t/instruction$3$_neg_lutinv }),
    .sr(rst_pad),
    .f({_al_u2802_o,open_n18373}),
    .q({open_n18377,\t/a/ID_op [3]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*A*(0@D))"),
    //.LUTF1("(0*~(C*~(~B*~(D*A))))"),
    //.LUTG0("(~C*~B*A*(1@D))"),
    //.LUTG1("(1*~(C*~(~B*~(D*A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b0001111100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2807|t/a/id_ex/reg5_b2  (
    .a({_al_u2801_o,_al_u2798_o}),
    .b({\t/a/n4_lutinv ,_al_u2799_o}),
    .c({\t/a/n2 ,_al_u2800_o}),
    .clk(clock_pad),
    .d({_al_u2806_o,_al_u2115_o}),
    .e({\t/busarbitration/n3_placeOpt_5 ,\t/a/ID_rd [2]}),
    .mi({open_n18380,\t/a/ID_rd [2]}),
    .sr(rst_pad),
    .f({_al_u2807_o,_al_u2801_o}),
    .q({open_n18395,\t/a/EX_rd [2]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("0"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111001111110011),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2808|t/a/id_ex/reg7_b9  (
    .b({open_n18398,\t/a/condition/n0_lutinv }),
    .c({open_n18399,\t/a/ID_memstraddr [9]}),
    .clk(clock_pad),
    .d({\t/a/condition/n0_lutinv ,\t/memstraddress [9]}),
    .e({_al_u2807_o,_al_u2807_o}),
    .mi({open_n18402,\t/a/ID_memstraddr [9]}),
    .sr(rst_pad),
    .f({_al_u2808_o,_al_u2812_o}),
    .q({open_n18417,\t/a/EX_memstraddr [9]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*D*~B*~C+A*D*~B*~C+~A*D*B*~C+A*D*B*~C"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~A*D*~B*~C+A*D*~B*~C+~A*D*B*~C+A*D*B*~C+~A*~D*~B*C+A*~D*~B*C+~A*D*~B*C+A*D*~B*C+~A*~D*B*C+A*~D*B*C+~A*D*B*C+A*D*B*C"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0111011101110111),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2809|t/a/if_id/reg5_b18  (
    .a({_al_u2792_o,open_n18418}),
    .b({_al_u2808_o,open_n18419}),
    .c({open_n18420,\t/busarbitration/n3_placeOpt_1 }),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({open_n18421,\t/a/MEM_aludat [18]}),
    .e({\t/instrnop ,\t/memstraddress [18]}),
    .mi({open_n18423,\t/memstraddress [18]}),
    .sr(rst_pad),
    .f({\t/a/if_id/n9 ,addr[18]}),
    .q({open_n18438,\t/a/ID_memstraddr [18]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("~B*~A*C*D+B*~A*C*D"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("~B*A*C*~D+B*A*C*~D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b0101000000000000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1111000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2811|_al_u2880  (
    .a({_al_u2810_o,n8[11]}),
    .b({open_n18439,_al_u2810_o}),
    .c({_al_u2109_o,\t/a/instr/n12 [12]}),
    .d({\t/a/instr/n16 [7],_al_u2109_o}),
    .e({n8[8],\t/a/instr/n16 [10]}),
    .f({_al_u2811_o,_al_u2880_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("D*B*C*~A+D*B*C*A"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("~D*~B*C*~A+D*~B*C*~A+D*B*C*~A+~D*~B*C*A+D*~B*C*A+D*B*C*A"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1111000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2814|_al_u2866  (
    .a({open_n18462,n8[16]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,\t/a/instr/n12 [17]}),
    .d({n8[7],_al_u2109_o}),
    .e({\t/a/instr/n16 [6],\t/a/instr/n16 [15]}),
    .f({_al_u2814_o,_al_u2866_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b1000100011110000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1011101111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2817|_al_u2854  (
    .a({n8[6],n8[20]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [7],\t/a/instr/n12 [21]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .e({\t/a/instr/n16 [5],\t/a/instr/n16 [19]}),
    .f({_al_u2817_o,_al_u2854_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b1000100011110000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1011101111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2819|_al_u2852  (
    .a({n8[5],n8[21]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [6],\t/a/instr/n12 [22]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .e({\t/a/instr/n16 [4],\t/a/instr/n16 [20]}),
    .f({_al_u2819_o,_al_u2852_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("A*B*C*~D+A*B*C*D"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b1000000010000000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1011000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2821|_al_u2831  (
    .a({n8[4],n8[2]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,\t/a/instr/n12 [3]}),
    .d({open_n18531,_al_u2109_o}),
    .e({\t/a/instr/n16 [3],\t/a/instr/n16 [1]}),
    .f({_al_u2821_o,_al_u2831_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b1000100011110000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1011101111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2824|_al_u2826  (
    .a({n8[3],n8[30]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [4],\t/a/instr/n12 [31]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .e({\t/a/instr/n16 [2],\t/a/instr/n16 [29]}),
    .f({_al_u2824_o,_al_u2826_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1011000010000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2828|_al_u2110  (
    .a({n8[29],_al_u2109_o}),
    .b({_al_u2810_o,\t/busarbitration/n3_placeOpt_4 }),
    .c({_al_u2109_o,\t/busarbitration/instruction [31]}),
    .clk(clock_pad),
    .d({\t/a/instr/n16 [28],i_data[31]}),
    .mi({i_data[31],i_data[31]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .f({_al_u2828_o,\t/a/IF_skip_addr [31]}),
    .q({\trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    //.LUT1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUT0(16'b1101000010000000),
    .INIT_LUT1(16'b1011000010000000),
    .MODE("LOGIC"))
    \_al_u2833|_al_u2887  (
    .a({n8[28],_al_u2810_o}),
    .b({_al_u2810_o,n8[0]}),
    .c({_al_u2109_o,_al_u2109_o}),
    .d({\t/a/instr/n16 [27],\t/memstraddress [1]}),
    .f({_al_u2833_o,_al_u2887_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUT1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUT0(16'b1000100011110000),
    .INIT_LUT1(16'b1011101111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2836 (
    .a({n8[27],n8[27]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [28],\t/a/instr/n12 [28]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .mi({open_n18620,\t/a/instr/n16 [26]}),
    .fx({open_n18625,_al_u2836_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUT1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUT0(16'b1000100011110000),
    .INIT_LUT1(16'b1011101111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2838 (
    .a({n8[26],n8[26]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [27],\t/a/instr/n12 [27]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .mi({open_n18640,\t/a/instr/n16 [25]}),
    .fx({open_n18645,_al_u2838_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1011000010000000),
    .MODE("LOGIC"))
    \_al_u2840|_al_u2810  (
    .a({n8[25],open_n18648}),
    .b({_al_u2810_o,open_n18649}),
    .c({_al_u2109_o,\t/a/condition/n0_lutinv }),
    .d({\t/a/instr/n16 [24],_al_u2792_o}),
    .f({_al_u2840_o,_al_u2810_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("A*D*B*~C+A*D*B*C"),
    //.LUTF1("D*A*B*~C+D*A*B*C"),
    //.LUTG0("~A*~D*B*~C+A*~D*B*~C+A*D*B*~C+~A*~D*B*C+A*~D*B*C+A*D*B*C"),
    //.LUTG1("~D*~A*B*~C+D*~A*B*~C+D*A*B*~C+~D*~A*B*C+D*~A*B*C+D*A*B*C"),
    .INIT_LUTF0(16'b1000100000000000),
    .INIT_LUTF1(16'b1000100000000000),
    .INIT_LUTG0(16'b1000100011001100),
    .INIT_LUTG1(16'b1100110001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2843|_al_u2882  (
    .a({_al_u2810_o,n8[10]}),
    .b({_al_u2109_o,_al_u2109_o}),
    .d({n8[24],_al_u2810_o}),
    .e({\t/a/instr/n16 [23],\t/a/instr/n16 [9]}),
    .f({_al_u2843_o,_al_u2882_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("D*B*C*~A+D*B*C*A"),
    //.LUTF1("~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG0("~D*~B*C*~A+D*~B*C*~A+D*B*C*~A+~D*~B*C*A+D*~B*C*A+D*B*C*A"),
    //.LUTG1("A*~C*B*~D+A*C*B*~D+A*~C*B*D+A*C*B*D"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100110000000000),
    .INIT_LUTG0(16'b1111000000110000),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2846|_al_u2877  (
    .a({n8[23],open_n18694}),
    .b({_al_u2109_o,_al_u2810_o}),
    .c({open_n18695,_al_u2109_o}),
    .d({\t/a/instr/n16 [22],n8[12]}),
    .e({_al_u2810_o,\t/a/instr/n16 [11]}),
    .f({_al_u2846_o,_al_u2877_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUT1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUT0(16'b1011000010000000),
    .INIT_LUT1(16'b1011000010000000),
    .MODE("LOGIC"))
    \_al_u2849|_al_u2874  (
    .a({n8[22],n8[13]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,_al_u2109_o}),
    .d({\t/a/instr/n16 [21],\t/a/instr/n16 [12]}),
    .f({_al_u2849_o,_al_u2874_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUT1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUT0(16'b1011000010000000),
    .INIT_LUT1(16'b1011000010000000),
    .MODE("LOGIC"))
    \_al_u2856|_al_u2871  (
    .a({n8[19],n8[14]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,_al_u2109_o}),
    .d({\t/a/instr/n16 [18],\t/a/instr/n16 [13]}),
    .f({_al_u2856_o,_al_u2871_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTF1("~A*~B*C*D+A*~B*C*D"),
    //.LUTG0("A*~B*C*~D+A*B*C*~D+A*~B*C*D+A*B*C*D"),
    //.LUTG1("~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b1010000010100000),
    .INIT_LUTG1(16'b1111000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2859|_al_u2868  (
    .a({open_n18758,n8[15]}),
    .b({_al_u2810_o,open_n18759}),
    .c({_al_u2109_o,_al_u2109_o}),
    .d({\t/a/instr/n16 [0],\t/a/instr/n16 [14]}),
    .e({n8[1],_al_u2810_o}),
    .f({_al_u2859_o,_al_u2868_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUT1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUT0(16'b1000100011110000),
    .INIT_LUT1(16'b1011101111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2862 (
    .a({n8[18],n8[18]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [19],\t/a/instr/n12 [19]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .mi({open_n18794,\t/a/instr/n16 [17]}),
    .fx({open_n18799,_al_u2862_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUT1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUT0(16'b1000100011110000),
    .INIT_LUT1(16'b1011101111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2864 (
    .a({n8[17],n8[17]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [18],\t/a/instr/n12 [18]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .mi({open_n18814,\t/a/instr/n16 [16]}),
    .fx({open_n18819,_al_u2864_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUT1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUT0(16'b1000100011110000),
    .INIT_LUT1(16'b1011101111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2885 (
    .a({n8[9],n8[9]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [10],\t/a/instr/n12 [10]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .mi({open_n18834,\t/a/instr/n16 [8]}),
    .fx({open_n18839,_al_u2885_o}));
  EG_PHY_GCLK _al_u2979 (
    .clki(jtck_leading),
    .clko(jtck));
  // D:/td/td/cw\register.v(31)
  EG_PHY_LSLICE #(
    //.LUTF0("C*~B*~A*D+C*B*~A*D+C*~B*A*D+C*B*A*D"),
    //.LUTF1("~A*B*D*~C+A*B*D*~C+~A*B*D*C+A*B*D*C"),
    //.LUTG0("~C*~B*~A*~D+~C*~B*A*~D+~C*~B*~A*D+C*~B*~A*D+C*B*~A*D+~C*~B*A*D+C*~B*A*D+C*B*A*D"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100110000000000),
    .INIT_LUTG0(16'b1111001100000011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3036|cfg_int/wrapper_cfg_inst/reg_inst/reg0_b17  (
    .b({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [0],_al_u3035_o}),
    .c({open_n18844,_al_u3034_o}),
    .clk(jtck),
    .d({_al_u3035_o,status_17}),
    .e({_al_u3034_o,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [17]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .f({jtdo_1,open_n18860}),
    .q({open_n18864,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [17]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_LSLICE #(
    //.LUTF0("0"),
    //.LUTF1("~A*~C*~D*~B+A*~C*~D*~B+~A*C*~D*~B+A*C*~D*~B+A*~C*D*~B+A*C*D*~B+~A*~C*~D*B+A*~C*~D*B+~A*C*~D*B+A*C*~D*B+A*~C*D*B+A*C*D*B"),
    //.LUTG0("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG1("~A*C*~D*~B+A*C*~D*~B+A*C*D*~B+~A*C*~D*B+A*C*~D*B+A*C*D*B"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010101011111111),
    .INIT_LUTG0(16'b1010101010101010),
    .INIT_LUTG1(16'b1010000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3057|_al_u3013  (
    .a({status_0,jshift}),
    .c({status_6,open_n18867}),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [0],open_n18870}),
    .e({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [6],jscan_0}),
    .f({_al_u3057_o,\cfg_int/wrapper_cfg_inst/shift_0 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*A)"),
    //.LUT1("(D*C*B*A)"),
    .INIT_LUT0(16'b0010001000100010),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"))
    \_al_u3062|_al_u3082  (
    .a({_al_u3056_o,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [12]}),
    .b({_al_u3058_o,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [12]}),
    .c({_al_u3060_o,open_n18891}),
    .d({_al_u3061_o,open_n18894}),
    .f({_al_u3062_o,_al_u3082_o}));
  // D:/td/td/cw\write_ctrl.v(36)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("~(~A*~B)"),
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3070|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/ce_reg  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n2 ,open_n18913}),
    .b({_al_u3069_o,open_n18914}),
    .c({open_n18915,\trig_node/trigger_node_int_0/pause_sync }),
    .clk(clock_pad),
    .d({open_n18917,status_17}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13$0$_en ,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n2 }),
    .q({open_n18933,wt_ce}));  // D:/td/td/cw\write_ctrl.v(36)
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~(~D*B)*~(C@A))"),
    //.LUTF1("~B*~C*~A*~D+~B*~C*A*~D+~B*~C*~A*D+~B*C*~A*D+~B*~C*A*D+~B*C*A*D"),
    //.LUTG0("(~1*~(~D*B)*~(C@A))"),
    //.LUTG1("~B*~C*~A*~D+B*~C*~A*~D+~B*~C*A*~D+B*~C*A*~D+~B*~C*~A*D+B*~C*~A*D+~B*C*~A*D+B*C*~A*D+~B*~C*A*D+B*~C*A*D+~B*C*A*D+B*C*A*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010010100100001),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3071|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b10  (
    .a({open_n18934,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [10]}),
    .b(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [10:9]),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [12],status_10}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [12],status_9}),
    .e({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [10],status_17}),
    .mi({open_n18937,status_10}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3071_o,_al_u3061_o}),
    .q({open_n18952,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [10]}));  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\write_ctrl.v(73)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~B)"),
    //.LUT1("(~D*A*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111011101110),
    .INIT_LUT1(16'b0000000010001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3072|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_reg  (
    .a({_al_u3071_o,status_17}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [2],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n19 }),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [2],open_n18953}),
    .clk(clock_pad),
    .d({status_17,open_n18955}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3072_o,open_n18968}),
    .q({open_n18972,status_17}));  // D:/td/td/cw\write_ctrl.v(73)
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*A)"),
    //.LUT1("(~(~D*B)*~(A*~C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3073|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b2  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [10],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [2]}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [2],open_n18973}),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [10],open_n18974}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [2],status_2}),
    .mi({open_n18986,status_2}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3073_o,_al_u3059_o}),
    .q({open_n18990,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [2]}));  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C@B)*~(D@A))"),
    //.LUT1("(B*C*~(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000001001000001),
    .INIT_LUT1(16'b1000000001000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3074|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b13  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [13],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [13]}),
    .b({_al_u3073_o,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [1]}),
    .c({_al_u3072_o,status_1}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [13],status_13}),
    .mi({open_n19002,status_13}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3074_o,_al_u3068_o}),
    .q({open_n19006,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [13]}));  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D@C)*~(~0*B))"),
    //.LUTF1("~B*A*~C*~D+B*A*~C*~D+~B*A*C*~D+B*A*C*~D"),
    //.LUTG0("(~A*~(D@C)*~(~1*B))"),
    //.LUTG1("~B*A*~C*D+B*A*~C*D+~B*A*C*D+B*A*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001000000000001),
    .INIT_LUTF1(16'b0000000010101010),
    .INIT_LUTG0(16'b0101000000000101),
    .INIT_LUTG1(16'b1010101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3076|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b4  (
    .a({_al_u3075_o,_al_u3059_o}),
    .b({open_n19007,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [8]}),
    .c({open_n19008,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [4]}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [4],status_4}),
    .e({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [4],status_8}),
    .mi({open_n19011,status_4}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3076_o,_al_u3060_o}),
    .q({open_n19026,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [4]}));  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~A)"),
    //.LUT1("(C*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010100000000),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3077|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b7  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [7],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [7]}),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [7],open_n19029}),
    .clk(clock_pad),
    .d({open_n19031,status_7}),
    .mi({open_n19042,status_7}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3077_o,_al_u3063_o}),
    .q({open_n19046,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [7]}));  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~C)*~(0*~B))"),
    //.LUTF1("~B*~A*~C*~D+~B*A*~C*~D+~B*A*~C*D"),
    //.LUTG0("(A*~(D*~C)*~(1*~B))"),
    //.LUTG1("~B*~A*C*~D+~B*A*C*~D+~B*A*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010000010101010),
    .INIT_LUTF1(16'b0000001000000011),
    .INIT_LUTG0(16'b1000000010001000),
    .INIT_LUTG1(16'b0010000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3078|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b8  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [8],_al_u3057_o}),
    .b({_al_u3077_o,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [8]}),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [0],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [2]}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [8],status_2}),
    .e({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [0],status_8}),
    .mi({open_n19049,status_8}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3078_o,_al_u3058_o}),
    .q({open_n19064,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [8]}));  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~B)*~(~D*A))"),
    //.LUT1("(~D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100111101000101),
    .INIT_LUT1(16'b0000000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3079|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b6  (
    .a({open_n19065,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [7]}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [6],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [6]}),
    .c({open_n19066,status_6}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [6],status_7}),
    .mi({open_n19078,status_6}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3079_o,_al_u3066_o}),
    .q({open_n19082,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [6]}));  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D@C)*~(~0*B))"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D+A*~C*B*~D+~A*C*~B*D+A*C*~B*D+A*C*B*D"),
    //.LUTG0("(~A*~(D@C)*~(~1*B))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001000000000001),
    .INIT_LUTF1(16'b1011000000001011),
    .INIT_LUTG0(16'b0101000000000101),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3080|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b11  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [7],_al_u3063_o}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [7],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [12]}),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [11],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [11]}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [11],status_11}),
    .e({_al_u3079_o,status_12}),
    .mi({open_n19085,status_11}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3080_o,_al_u3064_o}),
    .q({open_n19100,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [11]}));  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    .INIT_LUT0(16'b1000000000000000),
    .MODE("LOGIC"))
    _al_u3081 (
    .a({open_n19101,_al_u3074_o}),
    .b({open_n19102,_al_u3076_o}),
    .c({open_n19103,_al_u3078_o}),
    .d({open_n19106,_al_u3080_o}),
    .f({open_n19120,_al_u3081_o}));
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~A*~(D@C)*~(~0*B))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~A*~(D@C)*~(~1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0001000000000001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0101000000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3083|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b15  (
    .a({_al_u3082_o,_al_u3062_o}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [15],_al_u3067_o}),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [1],_al_u3068_o}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [1],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [15]}),
    .e({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [15],status_15}),
    .mi({open_n19128,status_15}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3083_o,_al_u3069_o}),
    .q({open_n19143,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [15]}));  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(A@C)*~(0*~B))"),
    //.LUTF1("0"),
    //.LUTG0("(~D*~(A@C)*~(1*~B))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D"),
    .INIT_LUTF0(16'b0000000010100101),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000010000100),
    .INIT_LUTG1(16'b0000000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u3084|_al_u3085  (
    .a({open_n19144,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [14]}),
    .b({open_n19145,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [15]}),
    .c({open_n19146,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [14]}),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [6],_al_u3084_o}),
    .e({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [6],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [15]}),
    .f({_al_u3084_o,_al_u3085_o}));
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~B)*~(D*~A))"),
    //.LUT1("(~(~A*B)*~(D@C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000101011001111),
    .INIT_LUT1(16'b1011000000001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3086|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b9  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [8],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [9]}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [8],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [0]}),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [9],status_0}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [9],status_9}),
    .mi({open_n19180,status_9}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3086_o,_al_u3055_o}),
    .q({open_n19184,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [9]}));  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("~C*B*A*D+C*B*A*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3120|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b93  (
    .a({_al_u3115_o,_al_u3108_o}),
    .b({_al_u3111_o,_al_u3109_o}),
    .c({open_n19185,_al_u3110_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3119_o,control_93}),
    .e({_al_u3107_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 }),
    .mi({open_n19187,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [93]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3120_o,_al_u3111_o}),
    .q({open_n19202,control_93}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(0*D*A*B*C)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(1*D*A*B*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3137|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b60  (
    .a({_al_u3128_o,_al_u3133_o}),
    .b({_al_u3124_o,_al_u3134_o}),
    .c({_al_u3120_o,_al_u3135_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3132_o,control_60}),
    .e({_al_u3136_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi({open_n19204,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [60]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3137_o,_al_u3136_o}),
    .q({open_n19219,control_60}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("A*B*C*D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3154|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b75  (
    .a({_al_u3141_o,_al_u3138_o}),
    .b({_al_u3153_o,_al_u3139_o}),
    .c({_al_u3145_o,_al_u3140_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3149_o,control_75}),
    .e({open_n19220,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi({open_n19222,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [75]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3154_o,_al_u3141_o}),
    .q({open_n19237,control_75}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(0*C*D*B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(1*C*D*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3171|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b276  (
    .a({_al_u3154_o,_al_u3155_o}),
    .b({_al_u3158_o,_al_u3156_o}),
    .c({_al_u3166_o,_al_u3157_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3162_o,control_276}),
    .e({_al_u3170_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi({open_n19239,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [276]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3171_o,_al_u3158_o}),
    .q({open_n19254,control_276}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("A*~D*C*B+A*D*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3188|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b90  (
    .a({_al_u3175_o,_al_u3172_o}),
    .b({_al_u3187_o,_al_u3173_o}),
    .c({_al_u3183_o,_al_u3174_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({open_n19255,control_90}),
    .e({_al_u3179_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 }),
    .mi({open_n19257,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [90]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3188_o,_al_u3175_o}),
    .q({open_n19272,control_90}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3197|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b72  (
    .a({_al_u3196_o,_al_u3189_o}),
    .b({_al_u3171_o,_al_u3190_o}),
    .c({_al_u3188_o,_al_u3191_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3192_o,control_72}),
    .e({_al_u3137_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({open_n19274,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [72]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3197_o,_al_u3192_o}),
    .q({open_n19289,control_72}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("D*C*A*~B+D*C*A*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3214|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b210  (
    .a({_al_u3209_o,_al_u3202_o}),
    .b({open_n19290,_al_u3203_o}),
    .c({_al_u3205_o,_al_u3204_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3201_o,control_210}),
    .e({_al_u3213_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({open_n19292,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [210]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3214_o,_al_u3205_o}),
    .q({open_n19307,control_210}));  // D:/td/td/cw\register.v(38)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1111001111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u322|_al_u1472  (
    .a({open_n19308,\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/busarbitration/n3_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/memstraddress [1],\t/a/regfile/regfile$0$ [1]}),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [1],\t/a/regfile/regfile$1$ [1]}),
    .mi({addr[1],addr[1]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .f({addr[1],_al_u1472_o}),
    .q({\trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/level_0_r }));
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3231|trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/ctl_last_reg  (
    .a({_al_u3214_o,control_211}),
    .b({_al_u3218_o,control_212}),
    .c({_al_u3222_o,\trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({_al_u3226_o,\trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/level_0_r }),
    .e({_al_u3230_o,\trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n19325,\trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .f({_al_u3231_o,_al_u3240_o}),
    .q({open_n19340,\trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUT1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111001001010000),
    .INIT_LUT1(16'b1111001111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u323|t/a/mem_wb/reg0_b0  (
    .a({open_n19341,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({\t/busarbitration/n3_placeOpt_2 ,_al_u1908_o}),
    .c({\t/memstraddress [0],\t/a/MEM_aludat [0]}),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [0],i_data[0]}),
    .sr(rst_pad),
    .f({addr[0],open_n19355}),
    .q({open_n19359,\t/a/reg_writedat [0]}));  // flow_line_reg.v(234)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("A*B*C*D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3248|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b216  (
    .a({_al_u3243_o,_al_u3244_o}),
    .b({_al_u3239_o,_al_u3245_o}),
    .c({_al_u3247_o,_al_u3246_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3235_o,control_216}),
    .e({open_n19360,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi({open_n19362,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [216]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .f({_al_u3248_o,_al_u3247_o}),
    .q({open_n19377,control_216}));  // D:/td/td/cw\register.v(38)
  EG_PHY_MSLICE #(
    //.LUT0("(C*A*D)"),
    //.LUT1("(A*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010000000000000),
    .INIT_LUT1(16'b1010000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u324|_al_u327  (
    .a({memwrite_cs,addr[2]}),
    .c({addr[5],memwrite_cs}),
    .clk(clock_pad),
    .d({n0,n0}),
    .mi({addr[5],addr[5]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .f({n2[3],n2[0]}),
    .q({\trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*A*B)"),
    //.LUT1("(A*C*B)"),
    .INIT_LUT0(16'b1000100000000000),
    .INIT_LUT1(16'b1000000010000000),
    .MODE("LOGIC"))
    \_al_u325|_al_u326  (
    .a({memwrite_cs,addr[3]}),
    .b({n0,n0}),
    .c({addr[4],open_n19394}),
    .d({open_n19397,memwrite_cs}),
    .f(n2[2:1]));
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(0*C*D*B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(1*C*D*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3265|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b27  (
    .a({_al_u3248_o,_al_u3257_o}),
    .b({_al_u3252_o,_al_u3258_o}),
    .c({_al_u3260_o,_al_u3259_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3256_o,control_27}),
    .e({_al_u3264_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({open_n19417,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [27]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3265_o,_al_u3260_o}),
    .q({open_n19432,control_27}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("D*A*C*~B+D*A*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3282|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b282  (
    .a({_al_u3273_o,_al_u3266_o}),
    .b({open_n19433,_al_u3267_o}),
    .c({_al_u3277_o,_al_u3268_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3269_o,control_282}),
    .e({_al_u3281_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi({open_n19435,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [282]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3282_o,_al_u3269_o}),
    .q({open_n19450,control_282}));  // D:/td/td/cw\register.v(38)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0@C)*~(D*~B))"),
    //.LUT1("(~A*~(1@B)*~(C*~D))"),
    .INIT_LUT0(16'b0000010000000101),
    .INIT_LUT1(16'b0100010000000100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u329 (
    .a({_al_u328_o,_al_u328_o}),
    .b({\t/a/ID_rs1 [3],\t/a/ID_rs1$0$_placeOpt_16 }),
    .c({\t/a/WB_rd [0],\t/a/ID_rs1 [3]}),
    .d({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/WB_rd [0]}),
    .mi({open_n19463,\t/a/WB_rd [3]}),
    .fx({open_n19468,_al_u329_o}));
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3299|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b87  (
    .a({_al_u3282_o,_al_u3295_o}),
    .b({_al_u3286_o,_al_u3296_o}),
    .c({_al_u3290_o,_al_u3297_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3294_o,control_87}),
    .e({_al_u3298_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({open_n19472,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [87]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3299_o,_al_u3298_o}),
    .q({open_n19487,control_87}));  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~C*~B*~A*~D+~C*B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*B*A*~D+C*B*A*~D+~C*~B*~A*D+~C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~C*~B*~A*D+~C*B*~A*D+~C*~B*A*D+C*~B*A*D+~C*B*A*D+C*B*A*D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1010111110101111),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1010111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u330|_al_u359  (
    .a({\t/a/WB_rd [0],_al_u355_o}),
    .b({open_n19488,_al_u356_o}),
    .c({\t/a/ID_rs1$0$_placeOpt_16 ,_al_u357_o}),
    .d({\t/a/WB_rd [4],_al_u358_o}),
    .e({\t/a/ID_rs1 [4],\t/a/ID_rs1$2$_placeOpt_9 }),
    .f({_al_u330_o,_al_u359_o}));
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("A*~B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3316|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b84  (
    .a({_al_u3303_o,_al_u3300_o}),
    .b({open_n19511,_al_u3301_o}),
    .c({_al_u3311_o,_al_u3302_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3315_o,control_84}),
    .e({_al_u3307_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({open_n19513,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [84]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3316_o,_al_u3303_o}),
    .q({open_n19528,control_84}));  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u331|_al_u915  (
    .a({\t/a/ID_rs1$1$_placeOpt_10 ,_al_u911_o}),
    .b({\t/a/ID_rs1 [4],_al_u912_o}),
    .c({\t/a/WB_rd [1],_al_u913_o}),
    .d({\t/a/WB_rd [4],_al_u914_o}),
    .e({open_n19531,\t/a/ID_rs1$2$_placeOpt_9 }),
    .f({_al_u331_o,_al_u915_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*A*~(0@D))"),
    //.LUT1("(C*B*A*~(1@D))"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u332 (
    .a({_al_u329_o,_al_u329_o}),
    .b({_al_u330_o,_al_u330_o}),
    .c({_al_u331_o,_al_u331_o}),
    .d({\t/a/ID_rs1$2$_placeOpt_6 ,\t/a/ID_rs1$2$_placeOpt_6 }),
    .mi({open_n19564,\t/a/WB_rd [2]}),
    .fx({open_n19569,\t/a/regfile/n1_lutinv }));
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(0*C*D*B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(1*C*D*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3333|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b51  (
    .a({_al_u3316_o,_al_u3321_o}),
    .b({_al_u3320_o,_al_u3322_o}),
    .c({_al_u3328_o,_al_u3323_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3324_o,control_51}),
    .e({_al_u3332_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi({open_n19573,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [51]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .f({_al_u3333_o,_al_u3324_o}),
    .q({open_n19588,control_51}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3334|trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/ctl_last_reg  (
    .a({_al_u3197_o,control_49}),
    .b({_al_u3231_o,control_50}),
    .c({_al_u3265_o,\trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({_al_u3299_o,\trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/level_0_r }),
    .e({_al_u3333_o,\trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n19591,\trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .f({_al_u3334_o,_al_u3321_o}),
    .q({open_n19606,\trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*~B*A)"),
    //.LUTF1("0"),
    //.LUTG0("(1*D*~C*~B*A)"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u333|_al_u2613  (
    .a({\t/a/regfile/n1_lutinv ,\t/a/regfile/n1_lutinv }),
    .b({open_n19607,\t/a/risk_jump/n24_lutinv }),
    .c({open_n19608,\t/a/risk_jump/n11_lutinv }),
    .d({open_n19611,\t/a/n19 }),
    .e({\t/a/WB_regwritecs ,\t/a/condition/n1_lutinv }),
    .f({_al_u333_o,_al_u2613_o}));
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("0"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("A*D*C*~B+A*D*C*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3351|trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/ctl_last_reg  (
    .a({_al_u3338_o,control_40}),
    .b({open_n19632,control_41}),
    .c({_al_u3346_o,\trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({_al_u3342_o,\trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/level_0_r }),
    .e({_al_u3350_o,\trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n19635,\trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .f({_al_u3351_o,_al_u3445_o}),
    .q({open_n19650,\trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3368|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b96  (
    .a({_al_u3351_o,_al_u3360_o}),
    .b({_al_u3355_o,_al_u3361_o}),
    .c({_al_u3359_o,_al_u3362_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3363_o,control_96}),
    .e({_al_u3367_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi({open_n19652,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [96]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3368_o,_al_u3363_o}),
    .q({open_n19667,control_96}));  // D:/td/td/cw\register.v(38)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u338 (
    .a({_al_u334_o,_al_u334_o}),
    .b({_al_u335_o,_al_u335_o}),
    .c({_al_u336_o,_al_u336_o}),
    .d({_al_u337_o,_al_u337_o}),
    .mi({open_n19680,\t/a/ID_rs1 [2]}),
    .fx({open_n19685,_al_u338_o}));
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("A*B*~C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3381|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b99  (
    .a({_al_u3368_o,_al_u3377_o}),
    .b({_al_u3372_o,_al_u3378_o}),
    .c({open_n19688,_al_u3379_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3380_o,control_99}),
    .e({_al_u3376_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi({open_n19690,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [99]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3381_o,_al_u3380_o}),
    .q({open_n19705,control_99}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("D*B*C*~A+D*B*C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3398|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b312  (
    .a({open_n19706,_al_u3390_o}),
    .b({_al_u3389_o,_al_u3391_o}),
    .c({_al_u3393_o,_al_u3392_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3385_o,control_312}),
    .e({_al_u3397_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi({open_n19708,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [312]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3398_o,_al_u3393_o}),
    .q({open_n19723,control_312}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(0*C*D*B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(1*C*D*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3415|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b309  (
    .a({_al_u3398_o,_al_u3403_o}),
    .b({_al_u3402_o,_al_u3404_o}),
    .c({_al_u3410_o,_al_u3405_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3406_o,control_309}),
    .e({_al_u3414_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi({open_n19725,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [309]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3415_o,_al_u3406_o}),
    .q({open_n19740,control_309}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("A*B*C*D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3432|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b45  (
    .a({_al_u3423_o,_al_u3428_o}),
    .b({_al_u3431_o,_al_u3429_o}),
    .c({_al_u3427_o,_al_u3430_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3419_o,control_45}),
    .e({open_n19741,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi({open_n19743,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [45]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3432_o,_al_u3431_o}),
    .q({open_n19758,control_45}));  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~A)*~(B)*~(D)+(~C*~A)*B*~(D)+~((~C*~A))*B*D+(~C*~A)*B*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~A)*~(B)*~(D)+(~C*~A)*B*~(D)+~((~C*~A))*B*D+(~C*~A)*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100110000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u343|t/a/regfile/reg0_b649  (
    .a({_al_u340_o,_al_u339_o}),
    .b({_al_u338_o,\t/a/ID_rs1$0$_placeOpt_7 }),
    .c({_al_u342_o,\t/a/ID_rs1$1$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$20$ [9]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [9]}),
    .mi({open_n19760,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u343_o,_al_u340_o}),
    .q({open_n19775,\t/a/regfile/regfile$20$ [9]}));  // register.v(63)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(0*C*D*B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(1*C*D*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3449|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b81  (
    .a({_al_u3432_o,_al_u3441_o}),
    .b({_al_u3436_o,_al_u3442_o}),
    .c({_al_u3444_o,_al_u3443_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3440_o,control_81}),
    .e({_al_u3448_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi({open_n19777,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [81]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3449_o,_al_u3444_o}),
    .q({open_n19792,control_81}));  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~D*~B*~A*~C+D*~B*~A*~C+~D*~B*A*~C+~D*~B*~A*C+D*~B*~A*C+~D*~B*A*C"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("D*~B*~A*~C+D*~B*~A*C"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0001000100110011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0001000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u344|_al_u411  (
    .a({\t/a/regfile/regfile$5$ [9],_al_u407_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_14 ,_al_u408_o}),
    .c({open_n19793,_al_u409_o}),
    .d({\t/a/ID_rs1$0$_placeOpt_14 ,_al_u410_o}),
    .e({\t/a/regfile/regfile$4$ [9],\t/a/ID_rs1$2$_placeOpt_7 }),
    .f({_al_u344_o,_al_u411_o}));
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("A*D*C*~B+A*D*C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3466|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b69  (
    .a({_al_u3453_o,_al_u3450_o}),
    .b({open_n19816,_al_u3451_o}),
    .c({_al_u3461_o,_al_u3452_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3457_o,control_69}),
    .e({_al_u3465_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi({open_n19818,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [69]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3466_o,_al_u3453_o}),
    .q({open_n19833,control_69}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(0*D*C*A*B)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(1*D*C*A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3483|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b255  (
    .a({_al_u3470_o,_al_u3479_o}),
    .b({_al_u3466_o,_al_u3480_o}),
    .c({_al_u3474_o,_al_u3481_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3478_o,control_255}),
    .e({_al_u3482_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi({open_n19835,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [255]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3483_o,_al_u3482_o}),
    .q({open_n19850,control_255}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("D*C*B*~A+D*C*B*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3500|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b273  (
    .a({open_n19851,_al_u3484_o}),
    .b({_al_u3495_o,_al_u3485_o}),
    .c({_al_u3491_o,_al_u3486_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3487_o,control_273}),
    .e({_al_u3499_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi({open_n19853,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [273]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3500_o,_al_u3487_o}),
    .q({open_n19868,control_273}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3517|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b294  (
    .a({_al_u3500_o,_al_u3513_o}),
    .b({_al_u3504_o,_al_u3514_o}),
    .c({_al_u3508_o,_al_u3515_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3512_o,control_294}),
    .e({_al_u3516_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi({open_n19870,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [294]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3517_o,_al_u3516_o}),
    .q({open_n19885,control_294}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3518|trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/ctl_last_reg  (
    .a({_al_u3381_o,control_307}),
    .b({_al_u3415_o,control_308}),
    .c({_al_u3449_o,\trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({_al_u3483_o,\trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/level_0_r }),
    .e({_al_u3517_o,\trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n19888,\trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .f({_al_u3518_o,_al_u3403_o}),
    .q({open_n19903,\trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~A*~B*~C*~D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("~A*~B*~C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3520|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b228  (
    .a({_al_u3201_o,_al_u3329_o}),
    .b({_al_u3205_o,_al_u3330_o}),
    .c({_al_u3209_o,_al_u3331_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3332_o,control_228}),
    .e({open_n19904,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({open_n19906,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [228]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3520_o,_al_u3332_o}),
    .q({open_n19921,control_228}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3521|trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/ctl_last_reg  (
    .a({_al_u3520_o,control_226}),
    .b({_al_u3218_o,control_227}),
    .c({_al_u3222_o,\trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({_al_u3226_o,\trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/level_0_r }),
    .e({_al_u3213_o,\trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n19924,\trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .f({_al_u3521_o,_al_u3329_o}),
    .q({open_n19939,\trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~A*~B*~C*~D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("~A*~B*~C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3522|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b213  (
    .a({_al_u3230_o,_al_u3240_o}),
    .b({_al_u3239_o,_al_u3241_o}),
    .c({_al_u3243_o,_al_u3242_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3235_o,control_213}),
    .e({open_n19940,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi({open_n19942,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [213]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .f({_al_u3522_o,_al_u3243_o}),
    .q({open_n19957,control_213}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~0*~D*~C*~A*B)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~1*~D*~C*~A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000100),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3523|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b231  (
    .a({_al_u3252_o,_al_u3249_o}),
    .b({_al_u3522_o,_al_u3250_o}),
    .c({_al_u3256_o,_al_u3251_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3260_o,control_231}),
    .e({_al_u3247_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({open_n19959,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [231]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3523_o,_al_u3252_o}),
    .q({open_n19974,control_231}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~C*~B*~A*~D+C*~B*~A*~D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000010001),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3524|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b264  (
    .a({_al_u3273_o,_al_u3270_o}),
    .b({_al_u3269_o,_al_u3271_o}),
    .c({open_n19975,_al_u3272_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3277_o,control_264}),
    .e({_al_u3170_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi({open_n19977,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [264]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3524_o,_al_u3273_o}),
    .q({open_n19992,control_264}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3525|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b78  (
    .a({_al_u3524_o,_al_u3291_o}),
    .b({_al_u3286_o,_al_u3292_o}),
    .c({_al_u3290_o,_al_u3293_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3294_o,control_78}),
    .e({_al_u3281_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi({open_n19994,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [78]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3525_o,_al_u3294_o}),
    .q({open_n20009,control_78}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~A*~B*~C*~D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("~A*~B*~C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3526|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b66  (
    .a({_al_u3307_o,_al_u3304_o}),
    .b({_al_u3303_o,_al_u3305_o}),
    .c({_al_u3298_o,_al_u3306_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3311_o,control_66}),
    .e({open_n20010,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({open_n20012,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [66]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3526_o,_al_u3307_o}),
    .q({open_n20027,control_66}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~0*~D*~C*~A*B)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~1*~D*~C*~A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000100),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3527|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b36  (
    .a({_al_u3320_o,_al_u3312_o}),
    .b({_al_u3526_o,_al_u3313_o}),
    .c({_al_u3324_o,_al_u3314_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3328_o,control_36}),
    .e({_al_u3315_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({open_n20029,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [36]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3527_o,_al_u3315_o}),
    .q({open_n20044,control_36}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3528|trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/ctl_last_reg  (
    .a({_al_u3521_o,control_229}),
    .b({_al_u3523_o,control_230}),
    .c({_al_u3525_o,\trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({_al_u3527_o,\trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/level_0_r }),
    .e({open_n20046,\trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n20048,\trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .f({_al_u3528_o,_al_u3249_o}),
    .q({open_n20063,\trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~B*~A*~C*~D+~B*A*~C*~D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3529|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b63  (
    .a({open_n20064,_al_u3176_o}),
    .b({_al_u3196_o,_al_u3177_o}),
    .c({_al_u3183_o,_al_u3178_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3179_o,control_63}),
    .e({_al_u3175_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({open_n20066,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [63]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3529_o,_al_u3179_o}),
    .q({open_n20081,control_63}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\trigger_node.v(82)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~A*~(C*B))"),
    //.LUT1("(~C*A)"),
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111101010),
    .INIT_LUT1(16'b0000101000001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3530|trig_node/trigger_node_int_0/emb_store_en_reg  (
    .a({_al_u3529_o,_al_u3519_o}),
    .b({open_n20082,_al_u3535_o}),
    .c({_al_u3192_o,_al_u3547_o}),
    .clk(clock_pad),
    .d({open_n20084,\trig_node/trigger_node_int_0/emb_store_en }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .f({_al_u3530_o,open_n20097}),
    .q({open_n20101,\trig_node/trigger_node_int_0/emb_store_en }));  // D:/td/td/cw\trigger_node.v(82)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~A*~D*~B*~C+~A*D*~B*~C"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000100000001),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3531|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b48  (
    .a({_al_u3187_o,_al_u3184_o}),
    .b({_al_u3111_o,_al_u3185_o}),
    .c({_al_u3115_o,_al_u3186_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({open_n20102,control_48}),
    .e({_al_u3107_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi({open_n20104,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [48]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3531_o,_al_u3187_o}),
    .q({open_n20119,control_48}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("0"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("~A*~B*~C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3532|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b54  (
    .a({_al_u3128_o,_al_u3116_o}),
    .b({_al_u3124_o,_al_u3117_o}),
    .c({_al_u3119_o,_al_u3118_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3132_o,control_54}),
    .e({_al_u3531_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi({open_n20121,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [54]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3532_o,_al_u3119_o}),
    .q({open_n20136,control_54}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~A*~B*~C*~D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("~A*~B*~C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3533|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b246  (
    .a({_al_u3145_o,_al_u3142_o}),
    .b({_al_u3141_o,_al_u3143_o}),
    .c({_al_u3136_o,_al_u3144_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3149_o,control_246}),
    .e({open_n20137,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi({open_n20139,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [246]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3533_o,_al_u3145_o}),
    .q({open_n20154,control_246}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~0*~D*~C*~A*B)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~1*~D*~C*~A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000100),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3534|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b249  (
    .a({_al_u3158_o,_al_u3163_o}),
    .b({_al_u3533_o,_al_u3164_o}),
    .c({_al_u3162_o,_al_u3165_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3166_o,control_249}),
    .e({_al_u3153_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi({open_n20156,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [249]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3534_o,_al_u3166_o}),
    .q({open_n20171,control_249}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("0"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3535|trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/ctl_last_reg  (
    .a({open_n20172,control_247}),
    .b({_al_u3530_o,control_248}),
    .c({_al_u3532_o,\trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({_al_u3534_o,\trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/level_0_r }),
    .e({_al_u3528_o,\trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n20175,\trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .f({_al_u3535_o,_al_u3163_o}),
    .q({open_n20190,\trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~A*~C*~D*~B+~A*~C*~D*B"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000101),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3536|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b42  (
    .a({_al_u3338_o,_al_u3445_o}),
    .b({open_n20191,_al_u3446_o}),
    .c({_al_u3342_o,_al_u3447_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3346_o,control_42}),
    .e({_al_u3448_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi({open_n20193,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [42]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3536_o,_al_u3448_o}),
    .q({open_n20208,control_42}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3537|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b219  (
    .a({_al_u3536_o,_al_u3356_o}),
    .b({_al_u3355_o,_al_u3357_o}),
    .c({_al_u3359_o,_al_u3358_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3363_o,control_219}),
    .e({_al_u3350_o,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi({open_n20210,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [219]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3537_o,_al_u3359_o}),
    .q({open_n20225,control_219}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3538|trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/ctl_last_reg  (
    .a({_al_u3537_o,control_217}),
    .b({_al_u3372_o,control_218}),
    .c({_al_u3376_o,\trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({_al_u3380_o,\trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/level_0_r }),
    .e({_al_u3367_o,\trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n20228,\trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .f({_al_u3538_o,_al_u3356_o}),
    .q({open_n20243,\trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~A*~D*~C*~B+~A*~D*~C*B"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000101),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3539|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b306  (
    .a({_al_u3385_o,_al_u3386_o}),
    .b({open_n20244,_al_u3387_o}),
    .c({_al_u3393_o,_al_u3388_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3389_o,control_306}),
    .e({_al_u3516_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi({open_n20246,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [306]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3539_o,_al_u3389_o}),
    .q({open_n20261,control_306}));  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000010111001100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u353|t/a/regfile/reg0_b393  (
    .a({_al_u350_o,_al_u349_o}),
    .b({_al_u348_o,\t/a/ID_rs1$0$_placeOpt_13 }),
    .c({_al_u352_o,\t/a/ID_rs1$1$_placeOpt_13 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$12$ [9]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [9]}),
    .mi({open_n20263,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u353_o,_al_u350_o}),
    .q({open_n20278,\t/a/regfile/regfile$12$ [9]}));  // register.v(63)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~0*~D*~C*~A*B)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~1*~D*~C*~A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000100),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3540|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b297  (
    .a({_al_u3402_o,_al_u3407_o}),
    .b({_al_u3539_o,_al_u3408_o}),
    .c({_al_u3406_o,_al_u3409_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3410_o,control_297}),
    .e({_al_u3397_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi({open_n20280,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [297]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3540_o,_al_u3410_o}),
    .q({open_n20295,control_297}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~A*~B*~C*~D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("~A*~B*~C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3541|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b300  (
    .a({_al_u3423_o,_al_u3411_o}),
    .b({_al_u3419_o,_al_u3412_o}),
    .c({_al_u3414_o,_al_u3413_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3427_o,control_300}),
    .e({open_n20296,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi({open_n20298,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [300]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3541_o,_al_u3414_o}),
    .q({open_n20313,control_300}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~0*~D*~C*~A*B)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~1*~D*~C*~A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000100),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3542|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b180  (
    .a({_al_u3436_o,_al_u3437_o}),
    .b({_al_u3541_o,_al_u3438_o}),
    .c({_al_u3440_o,_al_u3439_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3444_o,control_180}),
    .e({_al_u3431_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi({open_n20315,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [180]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3542_o,_al_u3440_o}),
    .q({open_n20330,control_180}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~B*~A*~C*~D+~B*~A*~C*D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000100000001),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3543|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b39  (
    .a({_al_u3457_o,_al_u3458_o}),
    .b({_al_u3453_o,_al_u3459_o}),
    .c({_al_u3461_o,_al_u3460_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({open_n20331,control_39}),
    .e({_al_u3264_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi({open_n20333,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [39]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3543_o,_al_u3461_o}),
    .q({open_n20348,control_39}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~0*~C*~D*~B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~1*~C*~D*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3544|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b57  (
    .a({_al_u3543_o,_al_u3462_o}),
    .b({_al_u3470_o,_al_u3463_o}),
    .c({_al_u3478_o,_al_u3464_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3474_o,control_57}),
    .e({_al_u3465_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi({open_n20350,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [57]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3544_o,_al_u3465_o}),
    .q({open_n20365,control_57}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3545|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b222  (
    .a({open_n20366,_al_u3492_o}),
    .b({_al_u3491_o,_al_u3493_o}),
    .c({_al_u3487_o,_al_u3494_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3495_o,control_222}),
    .e({_al_u3482_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi({open_n20368,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [222]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3545_o,_al_u3495_o}),
    .q({open_n20383,control_222}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \_al_u3546|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b288  (
    .a({_al_u3545_o,_al_u3505_o}),
    .b({_al_u3504_o,_al_u3506_o}),
    .c({_al_u3508_o,_al_u3507_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3512_o,control_288}),
    .e({_al_u3499_o,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi({open_n20385,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [288]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3546_o,_al_u3508_o}),
    .q({open_n20400,control_288}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u3547|trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/ctl_last_reg  (
    .a({_al_u3538_o,control_295}),
    .b({_al_u3540_o,control_296}),
    .c({_al_u3542_o,\trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({_al_u3544_o,\trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/level_0_r }),
    .e({_al_u3546_o,\trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n20403,\trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .f({_al_u3547_o,_al_u3407_o}),
    .q({open_n20418,\trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~D*~B*~A*~C+D*~B*~A*~C+~D*~B*A*~C+D*~B*A*~C+D*~B*~A*C+D*~B*A*C"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~D*~B*~A*~C+~D*~B*A*~C"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u355|_al_u1085  (
    .a({open_n20419,_al_u1081_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_15 ,_al_u1082_o}),
    .c({\t/a/regfile/regfile$4$ [8],_al_u1083_o}),
    .d({\t/a/ID_rs1$0$_placeOpt_15 ,_al_u1084_o}),
    .e({\t/a/regfile/regfile$5$ [8],\t/a/ID_rs2$2$_placeOpt_6 }),
    .f({_al_u355_o,_al_u1085_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u364|t/a/regfile/reg0_b392  (
    .a({_al_u359_o,_al_u360_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$0$_placeOpt_12 }),
    .c({_al_u363_o,\t/a/ID_rs1$1$_placeOpt_12 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u361_o,\t/a/regfile/regfile$12$ [8]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [8]}),
    .mi({open_n20443,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u364_o,_al_u361_o}),
    .q({open_n20458,\t/a/regfile/regfile$12$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u369|_al_u684  (
    .a({_al_u365_o,_al_u680_o}),
    .b({_al_u366_o,_al_u681_o}),
    .c({_al_u367_o,_al_u682_o}),
    .d({_al_u368_o,_al_u683_o}),
    .e({\t/a/ID_rs1$2$_placeOpt_7 ,\t/a/ID_rs1$2$_placeOpt_7 }),
    .f({_al_u369_o,_al_u684_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u374|t/a/regfile/reg0_b904  (
    .a({_al_u369_o,_al_u370_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_3 }),
    .c({_al_u373_o,\t/a/ID_rs1$1$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u371_o,\t/a/regfile/regfile$28$ [8]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [8]}),
    .mi({open_n20482,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u374_o,_al_u371_o}),
    .q({open_n20497,\t/a/regfile/regfile$28$ [8]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u380 (
    .a({_al_u376_o,_al_u376_o}),
    .b({_al_u377_o,_al_u377_o}),
    .c({_al_u378_o,_al_u378_o}),
    .d({_al_u379_o,_al_u379_o}),
    .mi({open_n20510,\t/a/ID_rs1 [2]}),
    .fx({open_n20515,_al_u380_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~A)*~(B)*~(D)+(~C*~A)*B*~(D)+~((~C*~A))*B*D+(~C*~A)*B*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~A)*~(B)*~(D)+(~C*~A)*B*~(D)+~((~C*~A))*B*D+(~C*~A)*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100110000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u385|t/a/regfile/reg0_b647  (
    .a({_al_u382_o,_al_u381_o}),
    .b({_al_u380_o,\t/a/ID_rs1$0$_placeOpt_7 }),
    .c({_al_u384_o,\t/a/ID_rs1$1$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$20$ [7]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [7]}),
    .mi({open_n20519,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({_al_u385_o,_al_u382_o}),
    .q({open_n20534,\t/a/regfile/regfile$20$ [7]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*D*~A*~C+B*D*~A*~C+B*D*A*~C+~B*D*~A*C+B*D*~A*C+B*D*A*C"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*A*C*~D+B*A*C*~D+~B*~A*~C*D+B*~A*~C*D"),
    //.LUTG0("~B*D*~A*~C+~B*D*~A*C"),
    //.LUTG1("0"),
    .INIT_LUTF0(16'b1101110100000000),
    .INIT_LUTF1(16'b0000010110101111),
    .INIT_LUTG0(16'b0001000100000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u386|_al_u1093  (
    .a({\t/a/ID_rs1$0$_placeOpt_1 ,\t/a/regfile/regfile$6$ [7]}),
    .b({open_n20535,\t/a/ID_rs2$0$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$4$ [7],open_n20536}),
    .d({\t/a/regfile/regfile$5$ [7],\t/a/ID_rs2$1$_placeOpt_13 }),
    .e({\t/a/ID_rs1$1$_placeOpt_1 ,\t/a/regfile/regfile$7$ [7]}),
    .f({_al_u386_o,_al_u1093_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u390 (
    .a({_al_u386_o,_al_u386_o}),
    .b({_al_u387_o,_al_u387_o}),
    .c({_al_u388_o,_al_u388_o}),
    .d({_al_u389_o,_al_u389_o}),
    .mi({open_n20571,\t/a/ID_rs1 [2]}),
    .fx({open_n20576,_al_u390_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000101000111010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u395|t/a/regfile/reg0_b391  (
    .a({_al_u390_o,_al_u391_o}),
    .b({_al_u394_o,\t/a/ID_rs1$0$_placeOpt_1 }),
    .c({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u392_o,\t/a/regfile/regfile$12$ [7]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [7]}),
    .mi({open_n20580,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({_al_u395_o,_al_u392_o}),
    .q({open_n20595,\t/a/regfile/regfile$12$ [7]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~A*~C)*~((~B*~D))*~(0)+(~A*~C)*(~B*~D)*~(0)+~((~A*~C))*(~B*~D)*0+(~A*~C)*(~B*~D)*0)"),
    //.LUTF1("~B*~C*~A*~D+B*~C*~A*~D+~B*C*~A*~D+~B*~C*A*~D+B*~C*A*~D+~B*C*A*~D"),
    //.LUTG0("~((~A*~C)*~((~B*~D))*~(1)+(~A*~C)*(~B*~D)*~(1)+~((~A*~C))*(~B*~D)*1+(~A*~C)*(~B*~D)*1)"),
    //.LUTG1("B*~C*~A*~D+B*~C*A*~D"),
    .INIT_LUTF0(16'b1111101011111010),
    .INIT_LUTF1(16'b0000000000111111),
    .INIT_LUTG0(16'b1111111111001100),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u397|_al_u401  (
    .a({open_n20596,_al_u400_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_18 ,_al_u398_o}),
    .c({\t/a/regfile/regfile$5$ [6],_al_u399_o}),
    .d({\t/a/ID_rs1$1$_placeOpt_18 ,_al_u397_o}),
    .e({\t/a/regfile/regfile$4$ [6],\t/a/ID_rs1$2$_placeOpt_3 }),
    .f({_al_u397_o,_al_u401_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u406|t/a/regfile/reg0_b390  (
    .a({_al_u401_o,_al_u402_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$0$_placeOpt_21 }),
    .c({_al_u405_o,\t/a/ID_rs1$1$_placeOpt_21 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u403_o,\t/a/regfile/regfile$12$ [6]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [6]}),
    .mi({open_n20620,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u406_o,_al_u403_o}),
    .q({open_n20635,\t/a/regfile/regfile$12$ [6]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u416|t/a/regfile/reg0_b902  (
    .a({_al_u411_o,_al_u412_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_15 }),
    .c({_al_u415_o,\t/a/ID_rs1$1$_placeOpt_15 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u413_o,\t/a/regfile/regfile$28$ [6]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [6]}),
    .mi({open_n20637,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u416_o,_al_u413_o}),
    .q({open_n20652,\t/a/regfile/regfile$28$ [6]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u422 (
    .a({_al_u418_o,_al_u418_o}),
    .b({_al_u419_o,_al_u419_o}),
    .c({_al_u420_o,_al_u420_o}),
    .d({_al_u421_o,_al_u421_o}),
    .mi({open_n20665,\t/a/ID_rs1$2$_placeOpt_9 }),
    .fx({open_n20670,_al_u422_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u427|t/a/regfile/reg0_b389  (
    .a({_al_u424_o,_al_u423_o}),
    .b({_al_u422_o,\t/a/ID_rs1$0$_placeOpt_18 }),
    .c({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$1$_placeOpt_18 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u426_o,\t/a/regfile/regfile$12$ [5]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [5]}),
    .mi({open_n20674,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u427_o,_al_u424_o}),
    .q({open_n20689,\t/a/regfile/regfile$12$ [5]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u432|_al_u621  (
    .a({_al_u428_o,_al_u617_o}),
    .b({_al_u429_o,_al_u618_o}),
    .c({_al_u430_o,_al_u619_o}),
    .d({_al_u431_o,_al_u620_o}),
    .e({\t/a/ID_rs1$2$_placeOpt_7 ,\t/a/ID_rs1$2$_placeOpt_7 }),
    .f({_al_u432_o,_al_u621_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u437|t/a/regfile/reg0_b901  (
    .a({_al_u434_o,_al_u433_o}),
    .b({_al_u432_o,\t/a/ID_rs1$0$_placeOpt_14 }),
    .c({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u436_o,\t/a/regfile/regfile$28$ [5]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [5]}),
    .mi({open_n20713,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u437_o,_al_u434_o}),
    .q({open_n20728,\t/a/regfile/regfile$28$ [5]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u443 (
    .a({_al_u439_o,_al_u439_o}),
    .b({_al_u440_o,_al_u440_o}),
    .c({_al_u441_o,_al_u441_o}),
    .d({_al_u442_o,_al_u442_o}),
    .mi({open_n20741,\t/a/ID_rs1 [2]}),
    .fx({open_n20746,_al_u443_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~A)*~(B)*~(D)+(~C*~A)*B*~(D)+~((~C*~A))*B*D+(~C*~A)*B*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~A)*~(B)*~(D)+(~C*~A)*B*~(D)+~((~C*~A))*B*D+(~C*~A)*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100110000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u448|t/a/regfile/reg0_b644  (
    .a({_al_u445_o,_al_u444_o}),
    .b({_al_u443_o,\t/a/ID_rs1$0$_placeOpt_5 }),
    .c({_al_u447_o,\t/a/ID_rs1$1$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$20$ [4]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [4]}),
    .mi({open_n20750,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u448_o,_al_u445_o}),
    .q({open_n20765,\t/a/regfile/regfile$20$ [4]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*~B*C*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*~C*D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0010001100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u449|_al_u453  (
    .a({\t/a/ID_rs1$0$_placeOpt_10 ,_al_u449_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_10 ,_al_u450_o}),
    .c({\t/a/regfile/regfile$4$ [4],_al_u451_o}),
    .d({open_n20768,_al_u452_o}),
    .e({\t/a/regfile/regfile$5$ [4],\t/a/ID_rs1$2$_placeOpt_9 }),
    .f({_al_u449_o,_al_u453_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+A*B*~C*D+A*B*C*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~A*B*~C*~D+~A*B*C*~D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1000100011001100),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000001000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u450|_al_u1159  (
    .a({\t/a/ID_rs1$0$_placeOpt_10 ,_al_u1155_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_10 ,_al_u1156_o}),
    .c({open_n20789,_al_u1157_o}),
    .d({\t/a/regfile/regfile$6$ [4],_al_u1158_o}),
    .e({\t/a/regfile/regfile$7$ [4],\t/a/ID_rs2$2$_placeOpt_10 }),
    .f({_al_u450_o,_al_u1159_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000010111001100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u458|t/a/regfile/reg0_b388  (
    .a({_al_u455_o,_al_u454_o}),
    .b({_al_u453_o,\t/a/ID_rs1$0$_placeOpt_13 }),
    .c({_al_u457_o,\t/a/ID_rs1$1$_placeOpt_13 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$12$ [4]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [4]}),
    .mi({open_n20813,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u458_o,_al_u455_o}),
    .q({open_n20828,\t/a/regfile/regfile$12$ [4]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~A*~C*~D*~B+A*~C*~D*~B+~A*~C*D*~B+A*~C*D*~B+~A*~C*~D*B+~A*~C*D*B"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("A*~C*~D*~B+A*~C*D*~B"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000011100000111),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000001000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u460|_al_u464  (
    .a({\t/a/ID_rs1$0$_placeOpt_1 ,_al_u460_o}),
    .b({\t/a/regfile/regfile$5$ [3],_al_u461_o}),
    .c({\t/a/ID_rs1$1$_placeOpt_1 ,_al_u462_o}),
    .d({open_n20831,_al_u463_o}),
    .e({\t/a/regfile/regfile$4$ [3],\t/a/ID_rs1$2$_placeOpt_9 }),
    .f({_al_u460_o,_al_u464_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000010111001100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u469|t/a/regfile/reg0_b387  (
    .a({_al_u466_o,_al_u465_o}),
    .b({_al_u464_o,\t/a/ID_rs1$0$_placeOpt_13 }),
    .c({_al_u468_o,\t/a/ID_rs1$1$_placeOpt_13 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$12$ [3]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [3]}),
    .mi({open_n20853,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u469_o,_al_u466_o}),
    .q({open_n20868,\t/a/regfile/regfile$12$ [3]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1101110111011000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1111111111111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u474|_al_u579  (
    .a({\t/a/ID_rs1 [2],_al_u575_o}),
    .b({_al_u471_o,_al_u576_o}),
    .c({_al_u472_o,_al_u577_o}),
    .d({_al_u473_o,_al_u578_o}),
    .e({_al_u470_o,\t/a/ID_rs1 [2]}),
    .f({_al_u474_o,_al_u579_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000010111001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u479|t/a/regfile/reg0_b899  (
    .a({_al_u476_o,_al_u475_o}),
    .b({_al_u474_o,\t/a/ID_rs1$0$_placeOpt_2 }),
    .c({_al_u478_o,\t/a/ID_rs1$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$28$ [3]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [3]}),
    .mi({open_n20892,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u479_o,_al_u476_o}),
    .q({open_n20907,\t/a/regfile/regfile$28$ [3]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u485 (
    .a({_al_u481_o,_al_u481_o}),
    .b({_al_u482_o,_al_u482_o}),
    .c({_al_u483_o,_al_u483_o}),
    .d({_al_u484_o,_al_u484_o}),
    .mi({open_n20920,\t/a/ID_rs1$2$_placeOpt_4 }),
    .fx({open_n20925,_al_u485_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~B*~D)*~(A)*~(C)+(~B*~D)*A*~(C)+~((~B*~D))*A*C+(~B*~D)*A*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~B*~D)*~(A)*~(C)+(~B*~D)*A*~(C)+~((~B*~D))*A*C+(~B*~D)*A*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010000010100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u490|t/a/regfile/reg0_b671  (
    .a({_al_u485_o,_al_u486_o}),
    .b({_al_u489_o,\t/a/ID_rs1$0$_placeOpt_10 }),
    .c({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u487_o,\t/a/regfile/regfile$20$ [31]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [31]}),
    .mi({open_n20929,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u490_o,_al_u487_o}),
    .q({open_n20944,\t/a/regfile/regfile$20$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u495 (
    .a({_al_u491_o,_al_u491_o}),
    .b({_al_u492_o,_al_u492_o}),
    .c({_al_u493_o,_al_u493_o}),
    .d({_al_u494_o,_al_u494_o}),
    .mi({open_n20957,\t/a/ID_rs1$2$_placeOpt_10 }),
    .fx({open_n20962,_al_u495_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000101000111010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u500|t/a/regfile/reg0_b415  (
    .a({_al_u495_o,_al_u496_o}),
    .b({_al_u499_o,\t/a/ID_rs1$0$_placeOpt_16 }),
    .c({\t/a/ID_rs1 [3],\t/a/ID_rs1$1$_placeOpt_16 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u497_o,\t/a/regfile/regfile$12$ [31]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [31]}),
    .mi({open_n20966,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u500_o,_al_u497_o}),
    .q({open_n20981,\t/a/regfile/regfile$12$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~D*~A*~C*~B+D*~A*~C*~B+~D*~A*~C*B+D*~A*~C*B"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~D*~A*~C*~B+D*~A*~C*~B+~D*~A*C*~B+D*~A*C*~B"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000010100000101),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0001000100010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u502|_al_u506  (
    .a({\t/a/ID_rs1$1$_placeOpt_20 ,_al_u502_o}),
    .b({\t/a/regfile/regfile$5$ [30],_al_u503_o}),
    .c({\t/a/regfile/regfile$4$ [30],_al_u504_o}),
    .d({open_n20984,_al_u505_o}),
    .e({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/ID_rs1$2$_placeOpt_9 }),
    .f({_al_u502_o,_al_u506_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000010111001100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u511|t/a/regfile/reg0_b414  (
    .a({_al_u508_o,_al_u507_o}),
    .b({_al_u506_o,\t/a/ID_rs1$0$_placeOpt_16 }),
    .c({_al_u510_o,\t/a/ID_rs1$1$_placeOpt_16 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [30]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [30]}),
    .mi({open_n21006,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u511_o,_al_u508_o}),
    .q({open_n21021,\t/a/regfile/regfile$12$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1011101110111000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1111111111111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u516|_al_u768  (
    .a({_al_u512_o,_al_u764_o}),
    .b({\t/a/ID_rs1 [2],_al_u765_o}),
    .c({_al_u514_o,_al_u766_o}),
    .d({_al_u515_o,_al_u767_o}),
    .e({_al_u513_o,\t/a/ID_rs1 [2]}),
    .f({_al_u516_o,_al_u768_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000101000111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u521|t/a/regfile/reg0_b926  (
    .a({_al_u516_o,_al_u517_o}),
    .b({_al_u520_o,\t/a/ID_rs1$0$_placeOpt_2 }),
    .c({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u518_o,\t/a/regfile/regfile$28$ [30]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [30]}),
    .mi({open_n21045,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u521_o,_al_u518_o}),
    .q({open_n21060,\t/a/regfile/regfile$28$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~A*~C)*~((~B*~D))*~(0)+(~A*~C)*(~B*~D)*~(0)+~((~A*~C))*(~B*~D)*0+(~A*~C)*(~B*~D)*0)"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D+~A*~C*B*~D+A*~C*B*~D+~A*~C*~B*D+~A*~C*B*D"),
    //.LUTG0("~((~A*~C)*~((~B*~D))*~(1)+(~A*~C)*(~B*~D)*~(1)+~((~A*~C))*(~B*~D)*1+(~A*~C)*(~B*~D)*1)"),
    //.LUTG1("A*~C*~B*~D+A*~C*B*~D"),
    .INIT_LUTF0(16'b1111101011111010),
    .INIT_LUTF1(16'b0000010100001111),
    .INIT_LUTG0(16'b1111111111001100),
    .INIT_LUTG1(16'b0000000000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u523|_al_u527  (
    .a({\t/a/ID_rs1$0$_placeOpt_10 ,_al_u526_o}),
    .b({open_n21061,_al_u524_o}),
    .c({\t/a/ID_rs1$1$_placeOpt_10 ,_al_u525_o}),
    .d({\t/a/regfile/regfile$5$ [2],_al_u523_o}),
    .e({\t/a/regfile/regfile$4$ [2],\t/a/ID_rs1$2$_placeOpt_9 }),
    .f({_al_u523_o,_al_u527_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u532|t/a/regfile/reg0_b386  (
    .a({_al_u527_o,_al_u528_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$0$_placeOpt_12 }),
    .c({_al_u531_o,\t/a/ID_rs1$1$_placeOpt_12 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u529_o,\t/a/regfile/regfile$12$ [2]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [2]}),
    .mi({open_n21085,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u532_o,_al_u529_o}),
    .q({open_n21100,\t/a/regfile/regfile$12$ [2]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u537 (
    .a({_al_u533_o,_al_u533_o}),
    .b({_al_u534_o,_al_u534_o}),
    .c({_al_u535_o,_al_u535_o}),
    .d({_al_u536_o,_al_u536_o}),
    .mi({open_n21113,\t/a/ID_rs1 [2]}),
    .fx({open_n21118,_al_u537_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000010111001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u542|t/a/regfile/reg0_b898  (
    .a({_al_u539_o,_al_u538_o}),
    .b({_al_u537_o,\t/a/ID_rs1$0$_placeOpt_19 }),
    .c({_al_u541_o,\t/a/ID_rs1$1$_placeOpt_19 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$28$ [2]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [2]}),
    .mi({open_n21122,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u542_o,_al_u539_o}),
    .q({open_n21137,\t/a/regfile/regfile$28$ [2]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u548 (
    .a({_al_u544_o,_al_u544_o}),
    .b({_al_u545_o,_al_u545_o}),
    .c({_al_u546_o,_al_u546_o}),
    .d({_al_u547_o,_al_u547_o}),
    .mi({open_n21150,\t/a/ID_rs1 [2]}),
    .fx({open_n21155,_al_u548_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~A)*~(B)*~(D)+(~C*~A)*B*~(D)+~((~C*~A))*B*D+(~C*~A)*B*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~A)*~(B)*~(D)+(~C*~A)*B*~(D)+~((~C*~A))*B*D+(~C*~A)*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100110000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u553|t/a/regfile/reg0_b669  (
    .a({_al_u550_o,_al_u549_o}),
    .b({_al_u548_o,\t/a/ID_rs1$0$_placeOpt_5 }),
    .c({_al_u552_o,\t/a/ID_rs1$1$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$20$ [29]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [29]}),
    .mi({open_n21159,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u553_o,_al_u550_o}),
    .q({open_n21174,\t/a/regfile/regfile$20$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*~B*C*D"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+D*~B*C*A"),
    //.LUTG0("~A*~B*~C*~D+~A*~B*~C*D"),
    //.LUTG1("~D*~B*~C*~A+~D*~B*~C*A"),
    .INIT_LUTF0(16'b0010001100100011),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0000000100000001),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u554|_al_u1260  (
    .a({open_n21175,\t/a/ID_rs2$0$_placeOpt_9 }),
    .b({\t/a/ID_rs1$1$_placeOpt_18 ,\t/a/ID_rs2$1$_placeOpt_18 }),
    .c({\t/a/regfile/regfile$4$ [29],\t/a/regfile/regfile$4$ [29]}),
    .d({\t/a/ID_rs1$0$_placeOpt_18 ,open_n21178}),
    .e({\t/a/regfile/regfile$5$ [29],\t/a/regfile/regfile$5$ [29]}),
    .f({_al_u554_o,_al_u1260_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u558|_al_u810  (
    .a({_al_u554_o,_al_u806_o}),
    .b({_al_u555_o,_al_u807_o}),
    .c({_al_u556_o,_al_u808_o}),
    .d({_al_u557_o,_al_u809_o}),
    .e({\t/a/ID_rs1$2$_placeOpt_3 ,\t/a/ID_rs1$2$_placeOpt_3 }),
    .f({_al_u558_o,_al_u810_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u563|t/a/regfile/reg0_b413  (
    .a({_al_u558_o,_al_u559_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$0$_placeOpt_12 }),
    .c({_al_u562_o,\t/a/ID_rs1$1$_placeOpt_12 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u560_o,\t/a/regfile/regfile$12$ [29]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [29]}),
    .mi({open_n21222,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u563_o,_al_u560_o}),
    .q({open_n21237,\t/a/regfile/regfile$12$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~A*~C)*~((~B*~D))*~(0)+(~A*~C)*(~B*~D)*~(0)+~((~A*~C))*(~B*~D)*0+(~A*~C)*(~B*~D)*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG0("~((~A*~C)*~((~B*~D))*~(1)+(~A*~C)*(~B*~D)*~(1)+~((~A*~C))*(~B*~D)*1+(~A*~C)*(~B*~D)*1)"),
    //.LUTG1("A*~B*~C*~D+A*~B*C*~D"),
    .INIT_LUTF0(16'b1111101011111010),
    .INIT_LUTF1(16'b0001000100110011),
    .INIT_LUTG0(16'b1111111111001100),
    .INIT_LUTG1(16'b0000000000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u565|_al_u569  (
    .a({\t/a/ID_rs1$0$_placeOpt_15 ,_al_u568_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_15 ,_al_u566_o}),
    .c({open_n21238,_al_u567_o}),
    .d({\t/a/regfile/regfile$5$ [28],_al_u565_o}),
    .e({\t/a/regfile/regfile$4$ [28],\t/a/ID_rs1$2$_placeOpt_1 }),
    .f({_al_u565_o,_al_u569_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000101000111010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u574|t/a/regfile/reg0_b412  (
    .a({_al_u569_o,_al_u570_o}),
    .b({_al_u573_o,\t/a/ID_rs1$0$_placeOpt_1 }),
    .c({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u571_o,\t/a/regfile/regfile$12$ [28]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [28]}),
    .mi({open_n21262,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u574_o,_al_u571_o}),
    .q({open_n21277,\t/a/regfile/regfile$12$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000010111001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u584|t/a/regfile/reg0_b924  (
    .a({_al_u581_o,_al_u580_o}),
    .b({_al_u579_o,\t/a/ID_rs1$0$_placeOpt_2 }),
    .c({_al_u583_o,\t/a/ID_rs1$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$28$ [28]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [28]}),
    .mi({open_n21279,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u584_o,_al_u581_o}),
    .q({open_n21294,\t/a/regfile/regfile$28$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u590|_al_u800  (
    .a({_al_u586_o,_al_u796_o}),
    .b({_al_u587_o,_al_u797_o}),
    .c({_al_u588_o,_al_u798_o}),
    .d({_al_u589_o,_al_u799_o}),
    .e({\t/a/ID_rs1$2$_placeOpt_2 ,\t/a/ID_rs1$2$_placeOpt_2 }),
    .f({_al_u590_o,_al_u800_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~A)*~(B)*~(D)+(~C*~A)*B*~(D)+~((~C*~A))*B*D+(~C*~A)*B*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~A)*~(B)*~(D)+(~C*~A)*B*~(D)+~((~C*~A))*B*D+(~C*~A)*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100110000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u595|t/a/regfile/reg0_b667  (
    .a({_al_u592_o,_al_u591_o}),
    .b({_al_u590_o,\t/a/ID_rs1$0$_placeOpt_7 }),
    .c({_al_u594_o,\t/a/ID_rs1$1$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$20$ [27]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [27]}),
    .mi({open_n21318,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u595_o,_al_u592_o}),
    .q({open_n21333,\t/a/regfile/regfile$20$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u600 (
    .a({_al_u596_o,_al_u596_o}),
    .b({_al_u597_o,_al_u597_o}),
    .c({_al_u598_o,_al_u598_o}),
    .d({_al_u599_o,_al_u599_o}),
    .mi({open_n21346,\t/a/ID_rs1$2$_placeOpt_9 }),
    .fx({open_n21351,_al_u600_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000010111001100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u605|t/a/regfile/reg0_b411  (
    .a({_al_u602_o,_al_u601_o}),
    .b({_al_u600_o,\t/a/ID_rs1$0$_placeOpt_13 }),
    .c({_al_u604_o,\t/a/ID_rs1$1$_placeOpt_13 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$12$ [27]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [27]}),
    .mi({open_n21355,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u605_o,_al_u602_o}),
    .q({open_n21370,\t/a/regfile/regfile$12$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*~B*~A*D+~C*~B*A*D"),
    //.LUTF1("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*~B*~A*D+~C*~B*A*D"),
    //.LUTG0("C*~B*~A*~D+C*~B*A*~D"),
    //.LUTG1("C*~B*~A*~D+C*~B*A*~D"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000000000110000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u607|_al_u1333  (
    .b({\t/a/ID_rs1$1$_placeOpt_18 ,\t/a/ID_rs2$1$_placeOpt_18 }),
    .c({\t/a/ID_rs1$0$_placeOpt_18 ,\t/a/ID_rs2$0$_placeOpt_20 }),
    .d({\t/a/regfile/regfile$5$ [26],\t/a/regfile/regfile$5$ [26]}),
    .e({\t/a/regfile/regfile$4$ [26],\t/a/regfile/regfile$4$ [26]}),
    .f({_al_u607_o,_al_u1333_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u611 (
    .a({_al_u607_o,_al_u607_o}),
    .b({_al_u608_o,_al_u608_o}),
    .c({_al_u609_o,_al_u609_o}),
    .d({_al_u610_o,_al_u610_o}),
    .mi({open_n21407,\t/a/ID_rs1$2$_placeOpt_8 }),
    .fx({open_n21412,_al_u611_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u616|t/a/regfile/reg0_b410  (
    .a({_al_u613_o,_al_u612_o}),
    .b({_al_u611_o,\t/a/ID_rs1$0$_placeOpt_9 }),
    .c({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u615_o,\t/a/regfile/regfile$12$ [26]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [26]}),
    .mi({open_n21416,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u616_o,_al_u613_o}),
    .q({open_n21431,\t/a/regfile/regfile$12$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u626|t/a/regfile/reg0_b922  (
    .a({_al_u623_o,_al_u622_o}),
    .b({_al_u621_o,\t/a/ID_rs1$0$_placeOpt_14 }),
    .c({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u625_o,\t/a/regfile/regfile$28$ [26]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [26]}),
    .mi({open_n21433,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u626_o,_al_u623_o}),
    .q({open_n21448,\t/a/regfile/regfile$28$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~A*~C)*~((~B*~D))*~(0)+(~A*~C)*(~B*~D)*~(0)+~((~A*~C))*(~B*~D)*0+(~A*~C)*(~B*~D)*0)"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D"),
    //.LUTG0("~((~A*~C)*~((~B*~D))*~(1)+(~A*~C)*(~B*~D)*~(1)+~((~A*~C))*(~B*~D)*1+(~A*~C)*(~B*~D)*1)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    .INIT_LUTF0(16'b1111101011111010),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b1111111111001100),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u628|_al_u632  (
    .a({\t/a/regfile/regfile$4$ [25],_al_u631_o}),
    .b({\t/a/regfile/regfile$5$ [25],_al_u629_o}),
    .c({open_n21449,_al_u630_o}),
    .d({\t/a/ID_rs1$1$_placeOpt_21 ,_al_u628_o}),
    .e({\t/a/ID_rs1$0$_placeOpt_21 ,\t/a/ID_rs1$2$_placeOpt_5 }),
    .f({_al_u628_o,_al_u632_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u637|t/a/regfile/reg0_b409  (
    .a({_al_u632_o,_al_u633_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$0$_placeOpt_21 }),
    .c({_al_u636_o,\t/a/ID_rs1$1$_placeOpt_21 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u634_o,\t/a/regfile/regfile$12$ [25]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [25]}),
    .mi({open_n21473,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u637_o,_al_u634_o}),
    .q({open_n21488,\t/a/regfile/regfile$12$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u642 (
    .a({_al_u638_o,_al_u638_o}),
    .b({_al_u639_o,_al_u639_o}),
    .c({_al_u640_o,_al_u640_o}),
    .d({_al_u641_o,_al_u641_o}),
    .mi({open_n21501,\t/a/ID_rs1$2$_placeOpt_5 }),
    .fx({open_n21506,_al_u642_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u647|t/a/regfile/reg0_b921  (
    .a({_al_u642_o,_al_u643_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_21 }),
    .c({_al_u646_o,\t/a/ID_rs1$1$_placeOpt_21 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u644_o,\t/a/regfile/regfile$28$ [25]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [25]}),
    .mi({open_n21510,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u647_o,_al_u644_o}),
    .q({open_n21525,\t/a/regfile/regfile$28$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u653|_al_u957  (
    .a({_al_u649_o,_al_u953_o}),
    .b({_al_u650_o,_al_u954_o}),
    .c({_al_u651_o,_al_u955_o}),
    .d({_al_u652_o,_al_u956_o}),
    .e({\t/a/ID_rs1$2$_placeOpt_5 ,\t/a/ID_rs1$2$_placeOpt_5 }),
    .f({_al_u653_o,_al_u957_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000101000111010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u658|t/a/regfile/reg0_b408  (
    .a({_al_u653_o,_al_u654_o}),
    .b({_al_u657_o,\t/a/ID_rs1$0$_placeOpt_1 }),
    .c({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u655_o,\t/a/regfile/regfile$12$ [24]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [24]}),
    .mi({open_n21549,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u658_o,_al_u655_o}),
    .q({open_n21564,\t/a/regfile/regfile$12$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u663 (
    .a({_al_u659_o,_al_u659_o}),
    .b({_al_u660_o,_al_u660_o}),
    .c({_al_u661_o,_al_u661_o}),
    .d({_al_u662_o,_al_u662_o}),
    .mi({open_n21577,\t/a/ID_rs1$2$_placeOpt_7 }),
    .fx({open_n21582,_al_u663_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u668|t/a/regfile/reg0_b920  (
    .a({_al_u663_o,_al_u664_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_14 }),
    .c({_al_u667_o,\t/a/ID_rs1$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u665_o,\t/a/regfile/regfile$28$ [24]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [24]}),
    .mi({open_n21586,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u668_o,_al_u665_o}),
    .q({open_n21601,\t/a/regfile/regfile$28$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~A*~C)*~((~B*~D))*~(0)+(~A*~C)*(~B*~D)*~(0)+~((~A*~C))*(~B*~D)*0+(~A*~C)*(~B*~D)*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    //.LUTG0("~((~A*~C)*~((~B*~D))*~(1)+(~A*~C)*(~B*~D)*~(1)+~((~A*~C))*(~B*~D)*1+(~A*~C)*(~B*~D)*1)"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*C*~D"),
    .INIT_LUTF0(16'b1111101011111010),
    .INIT_LUTF1(16'b0010001000110011),
    .INIT_LUTG0(16'b1111111111001100),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u670|_al_u674  (
    .a({\t/a/ID_rs1$0$_placeOpt_12 ,_al_u673_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_12 ,_al_u671_o}),
    .c({open_n21602,_al_u672_o}),
    .d({\t/a/regfile/regfile$4$ [23],_al_u670_o}),
    .e({\t/a/regfile/regfile$5$ [23],\t/a/ID_rs1$2$_placeOpt_8 }),
    .f({_al_u670_o,_al_u674_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u679|t/a/regfile/reg0_b407  (
    .a({_al_u676_o,_al_u675_o}),
    .b({_al_u674_o,\t/a/ID_rs1$0$_placeOpt_12 }),
    .c({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$1$_placeOpt_12 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u678_o,\t/a/regfile/regfile$12$ [23]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [23]}),
    .mi({open_n21626,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u679_o,_al_u676_o}),
    .q({open_n21641,\t/a/regfile/regfile$12$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u689|t/a/regfile/reg0_b919  (
    .a({_al_u684_o,_al_u685_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .c({_al_u688_o,\t/a/ID_rs1$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u686_o,\t/a/regfile/regfile$28$ [23]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [23]}),
    .mi({open_n21643,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u689_o,_al_u686_o}),
    .q({open_n21658,\t/a/regfile/regfile$28$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u695|_al_u947  (
    .a({_al_u691_o,_al_u943_o}),
    .b({_al_u692_o,_al_u944_o}),
    .c({_al_u693_o,_al_u945_o}),
    .d({_al_u694_o,_al_u946_o}),
    .e({\t/a/ID_rs1$2$_placeOpt_7 ,\t/a/ID_rs1$2$_placeOpt_7 }),
    .f({_al_u695_o,_al_u947_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~B*~D)*~(A)*~(C)+(~B*~D)*A*~(C)+~((~B*~D))*A*C+(~B*~D)*A*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~B*~D)*~(A)*~(C)+(~B*~D)*A*~(C)+~((~B*~D))*A*C+(~B*~D)*A*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010000010100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u700|t/a/regfile/reg0_b662  (
    .a({_al_u695_o,_al_u696_o}),
    .b({_al_u699_o,\t/a/ID_rs1$0$_placeOpt_8 }),
    .c({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u697_o,\t/a/regfile/regfile$20$ [22]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [22]}),
    .mi({open_n21682,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u700_o,_al_u697_o}),
    .q({open_n21697,\t/a/regfile/regfile$20$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000000000110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u701|t/a/regfile/reg0_b182  (
    .a({\t/a/regfile/regfile$4$ [22],_al_u1853_o}),
    .b({\t/a/regfile/regfile$5$ [22],\t/a/alu_A_select [1]}),
    .c({\t/a/ID_rs1$0$_placeOpt_15 ,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_15 ,\t/a/reg_writedat [22]}),
    .mi({open_n21708,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u701_o,\t/a/aluin/sel0_b22/B0 }),
    .q({open_n21712,\t/a/regfile/regfile$5$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1101110111011000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1111111111111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u705|_al_u1411  (
    .a({\t/a/ID_rs1$2$_placeOpt_1 ,_al_u1407_o}),
    .b({_al_u702_o,_al_u1408_o}),
    .c({_al_u703_o,_al_u1409_o}),
    .d({_al_u704_o,_al_u1410_o}),
    .e({_al_u701_o,\t/a/ID_rs2$2$_placeOpt_6 }),
    .f({_al_u705_o,_al_u1411_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~C*~A))*~(D)+B*(~C*~A)*~(D)+~(B)*(~C*~A)*D+B*(~C*~A)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000010111001100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u710|t/a/regfile/reg0_b406  (
    .a({_al_u707_o,_al_u706_o}),
    .b({_al_u705_o,\t/a/ID_rs1$0$_placeOpt_13 }),
    .c({_al_u709_o,\t/a/ID_rs1$1$_placeOpt_13 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/regfile/regfile$12$ [22]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [22]}),
    .mi({open_n21736,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u710_o,_al_u707_o}),
    .q({open_n21751,\t/a/regfile/regfile$12$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u712|t/a/regfile/reg0_b181  (
    .a({\t/a/ID_rs1$0$_placeOpt_15 ,_al_u1856_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_15 ,\t/a/alu_A_select [1]}),
    .c({\t/a/regfile/regfile$4$ [21],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [21],\t/a/reg_writedat [21]}),
    .mi({open_n21762,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u712_o,\t/a/aluin/sel0_b21/B0 }),
    .q({open_n21766,\t/a/regfile/regfile$5$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u716 (
    .a({_al_u712_o,_al_u712_o}),
    .b({_al_u713_o,_al_u713_o}),
    .c({_al_u714_o,_al_u714_o}),
    .d({_al_u715_o,_al_u715_o}),
    .mi({open_n21779,\t/a/ID_rs1$2$_placeOpt_5 }),
    .fx({open_n21784,_al_u716_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u721|t/a/regfile/reg0_b405  (
    .a({_al_u716_o,_al_u717_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .c({_al_u720_o,\t/a/ID_rs1$1$_placeOpt_11 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u718_o,\t/a/regfile/regfile$12$ [21]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [21]}),
    .mi({open_n21788,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u721_o,_al_u718_o}),
    .q({open_n21803,\t/a/regfile/regfile$12$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u726 (
    .a({_al_u722_o,_al_u722_o}),
    .b({_al_u723_o,_al_u723_o}),
    .c({_al_u724_o,_al_u724_o}),
    .d({_al_u725_o,_al_u725_o}),
    .mi({open_n21816,\t/a/ID_rs1$2$_placeOpt_7 }),
    .fx({open_n21821,_al_u726_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u731|t/a/regfile/reg0_b917  (
    .a({_al_u726_o,_al_u727_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .c({_al_u730_o,\t/a/ID_rs1$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u728_o,\t/a/regfile/regfile$28$ [21]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [21]}),
    .mi({open_n21825,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u731_o,_al_u728_o}),
    .q({open_n21840,\t/a/regfile/regfile$28$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u737|_al_u905  (
    .a({_al_u733_o,_al_u901_o}),
    .b({_al_u734_o,_al_u902_o}),
    .c({_al_u735_o,_al_u903_o}),
    .d({_al_u736_o,_al_u904_o}),
    .e({\t/a/ID_rs1$2$_placeOpt_2 ,\t/a/ID_rs1$2$_placeOpt_2 }),
    .f({_al_u737_o,_al_u905_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~B*~D)*~(A)*~(C)+(~B*~D)*A*~(C)+~((~B*~D))*A*C+(~B*~D)*A*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~B*~D)*~(A)*~(C)+(~B*~D)*A*~(C)+~((~B*~D))*A*C+(~B*~D)*A*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010000010100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u742|t/a/regfile/reg0_b660  (
    .a({_al_u737_o,_al_u738_o}),
    .b({_al_u741_o,\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u739_o,\t/a/regfile/regfile$20$ [20]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [20]}),
    .mi({open_n21864,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u742_o,_al_u739_o}),
    .q({open_n21879,\t/a/regfile/regfile$20$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u747|_al_u863  (
    .a({_al_u743_o,_al_u859_o}),
    .b({_al_u744_o,_al_u860_o}),
    .c({_al_u745_o,_al_u861_o}),
    .d({_al_u746_o,_al_u862_o}),
    .e({\t/a/ID_rs1$2$_placeOpt_3 ,\t/a/ID_rs1$2$_placeOpt_3 }),
    .f({_al_u747_o,_al_u863_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u752|t/a/regfile/reg0_b404  (
    .a({_al_u747_o,_al_u748_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$0$_placeOpt_18 }),
    .c({_al_u751_o,\t/a/ID_rs1$1$_placeOpt_18 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u749_o,\t/a/regfile/regfile$12$ [20]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [20]}),
    .mi({open_n21903,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u752_o,_al_u749_o}),
    .q({open_n21918,\t/a/regfile/regfile$12$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~B*~D*~A*~C+B*~D*~A*~C+B*~D*A*~C+~B*~D*~A*C+B*~D*~A*C+B*~D*A*C"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~B*~D*~A*~C+~B*~D*~A*C"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000011011101),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u754|_al_u758  (
    .a({\t/a/regfile/regfile$4$ [1],_al_u754_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_16 ,_al_u755_o}),
    .c({open_n21919,_al_u756_o}),
    .d({\t/a/ID_rs1$1$_placeOpt_16 ,_al_u757_o}),
    .e({\t/a/regfile/regfile$5$ [1],\t/a/ID_rs1$2$_placeOpt_6 }),
    .f({_al_u754_o,_al_u758_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000101000111010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u763|t/a/regfile/reg0_b385  (
    .a({_al_u758_o,_al_u759_o}),
    .b({_al_u762_o,\t/a/ID_rs1$0$_placeOpt_16 }),
    .c({\t/a/ID_rs1 [3],\t/a/ID_rs1$1$_placeOpt_16 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u760_o,\t/a/regfile/regfile$12$ [1]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [1]}),
    .mi({open_n21943,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u763_o,_al_u760_o}),
    .q({open_n21958,\t/a/regfile/regfile$12$ [1]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~B*~D))*~(C)+A*(~B*~D)*~(C)+~(A)*(~B*~D)*C+A*(~B*~D)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000101000111010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u773|t/a/regfile/reg0_b897  (
    .a({_al_u768_o,_al_u769_o}),
    .b({_al_u772_o,\t/a/ID_rs1$0$_placeOpt_19 }),
    .c({\t/a/ID_rs1$3$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_19 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u770_o,\t/a/regfile/regfile$28$ [1]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [1]}),
    .mi({open_n21960,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u773_o,_al_u770_o}),
    .q({open_n21975,\t/a/regfile/regfile$28$ [1]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*C*~D+~A*B*C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTF1("~C*~B*~D*~A+C*~B*~D*~A+~C*~B*D*~A+~C*~B*~D*A+C*~B*~D*A+~C*~B*D*A"),
    //.LUTG0("~A*~B*C*D+~A*B*C*D"),
    //.LUTG1("C*~B*~D*~A+C*~B*~D*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000001010000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0101000000000000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u775|t/a/regfile/reg0_b179  (
    .a({open_n21976,_al_u1865_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_15 ,open_n21977}),
    .c({\t/a/ID_rs1$0$_placeOpt_15 ,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [19],\t/a/reg_writedat [19]}),
    .e({\t/a/regfile/regfile$4$ [19],\t/a/alu_A_select [1]}),
    .mi({open_n21979,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u775_o,\t/a/aluin/sel0_b19/B0 }),
    .q({open_n21994,\t/a/regfile/regfile$5$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u779 (
    .a({_al_u775_o,_al_u775_o}),
    .b({_al_u776_o,_al_u776_o}),
    .c({_al_u777_o,_al_u777_o}),
    .d({_al_u778_o,_al_u778_o}),
    .mi({open_n22007,\t/a/ID_rs1$2$_placeOpt_3 }),
    .fx({open_n22012,_al_u779_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u784|t/a/regfile/reg0_b403  (
    .a({_al_u779_o,_al_u780_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .c({_al_u783_o,\t/a/ID_rs1$1$_placeOpt_17 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u781_o,\t/a/regfile/regfile$12$ [19]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [19]}),
    .mi({open_n22016,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u784_o,_al_u781_o}),
    .q({open_n22031,\t/a/regfile/regfile$12$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u789 (
    .a({_al_u785_o,_al_u785_o}),
    .b({_al_u786_o,_al_u786_o}),
    .c({_al_u787_o,_al_u787_o}),
    .d({_al_u788_o,_al_u788_o}),
    .mi({open_n22044,\t/a/ID_rs1$2$_placeOpt_7 }),
    .fx({open_n22049,_al_u789_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u794|t/a/regfile/reg0_b915  (
    .a({_al_u791_o,_al_u790_o}),
    .b({_al_u789_o,\t/a/ID_rs1$0$_placeOpt_14 }),
    .c({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u793_o,\t/a/regfile/regfile$28$ [19]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [19]}),
    .mi({open_n22053,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u794_o,_al_u791_o}),
    .q({open_n22068,\t/a/regfile/regfile$28$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100000011000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u805|t/a/regfile/reg0_b658  (
    .a({_al_u802_o,_al_u801_o}),
    .b({_al_u800_o,\t/a/ID_rs1$0$_placeOpt_6 }),
    .c({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u804_o,\t/a/regfile/regfile$20$ [18]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [18]}),
    .mi({open_n22070,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u805_o,_al_u802_o}),
    .q({open_n22085,\t/a/regfile/regfile$20$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u806|t/a/regfile/reg0_b178  (
    .a({\t/a/regfile/regfile$5$ [18],_al_u1868_o}),
    .b({\t/a/regfile/regfile$4$ [18],\t/a/alu_A_select [1]}),
    .c({\t/a/ID_rs1$1$_placeOpt_15 ,\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_15 ,\t/a/reg_writedat [18]}),
    .mi({open_n22096,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u806_o,\t/a/aluin/sel0_b18/B0 }),
    .q({open_n22100,\t/a/regfile/regfile$5$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u815|t/a/regfile/reg0_b402  (
    .a({_al_u810_o,_al_u811_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$0$_placeOpt_21 }),
    .c({_al_u814_o,\t/a/ID_rs1$1$_placeOpt_21 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u812_o,\t/a/regfile/regfile$12$ [18]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [18]}),
    .mi({open_n22102,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u815_o,_al_u812_o}),
    .q({open_n22117,\t/a/regfile/regfile$12$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u821 (
    .a({_al_u817_o,_al_u817_o}),
    .b({_al_u818_o,_al_u818_o}),
    .c({_al_u819_o,_al_u819_o}),
    .d({_al_u820_o,_al_u820_o}),
    .mi({open_n22130,\t/a/ID_rs1$2$_placeOpt_5 }),
    .fx({open_n22135,_al_u821_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u826|t/a/regfile/reg0_b401  (
    .a({_al_u823_o,_al_u822_o}),
    .b({_al_u821_o,\t/a/ID_rs1$0$_placeOpt_11 }),
    .c({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u825_o,\t/a/regfile/regfile$12$ [17]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [17]}),
    .mi({open_n22139,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u826_o,_al_u823_o}),
    .q({open_n22154,\t/a/regfile/regfile$12$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u831|_al_u873  (
    .a({_al_u827_o,_al_u869_o}),
    .b({_al_u828_o,_al_u870_o}),
    .c({_al_u829_o,_al_u871_o}),
    .d({_al_u830_o,_al_u872_o}),
    .e({\t/a/ID_rs1$2$_placeOpt_5 ,\t/a/ID_rs1$2$_placeOpt_5 }),
    .f({_al_u831_o,_al_u873_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u836|t/a/regfile/reg0_b913  (
    .a({_al_u833_o,_al_u832_o}),
    .b({_al_u831_o,\t/a/ID_rs1$0$_placeOpt_14 }),
    .c({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u835_o,\t/a/regfile/regfile$28$ [17]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [17]}),
    .mi({open_n22178,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u836_o,_al_u833_o}),
    .q({open_n22193,\t/a/regfile/regfile$28$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u842 (
    .a({_al_u838_o,_al_u838_o}),
    .b({_al_u839_o,_al_u839_o}),
    .c({_al_u840_o,_al_u840_o}),
    .d({_al_u841_o,_al_u841_o}),
    .mi({open_n22206,\t/a/ID_rs1$2$_placeOpt_2 }),
    .fx({open_n22211,_al_u842_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~D*~A)*~(B)*~(C)+(~D*~A)*B*~(C)+~((~D*~A))*B*C+(~D*~A)*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100000011000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u847|t/a/regfile/reg0_b656  (
    .a({_al_u844_o,_al_u843_o}),
    .b({_al_u842_o,\t/a/ID_rs1$0$_placeOpt_3 }),
    .c({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u846_o,\t/a/regfile/regfile$20$ [16]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [16]}),
    .mi({open_n22215,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u847_o,_al_u844_o}),
    .q({open_n22230,\t/a/regfile/regfile$20$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u852|_al_u1558  (
    .a({_al_u848_o,_al_u1554_o}),
    .b({_al_u849_o,_al_u1555_o}),
    .c({_al_u850_o,_al_u1556_o}),
    .d({_al_u851_o,_al_u1557_o}),
    .e({\t/a/ID_rs1$2$_placeOpt_3 ,\t/a/ID_rs2$2$_placeOpt_3 }),
    .f({_al_u852_o,_al_u1558_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u857|t/a/regfile/reg0_b400  (
    .a({_al_u854_o,_al_u853_o}),
    .b({_al_u852_o,\t/a/ID_rs1$0$_placeOpt_18 }),
    .c({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$1$_placeOpt_18 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u856_o,\t/a/regfile/regfile$12$ [16]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [16]}),
    .mi({open_n22254,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u857_o,_al_u854_o}),
    .q({open_n22269,\t/a/regfile/regfile$12$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u868|t/a/regfile/reg0_b399  (
    .a({_al_u865_o,_al_u864_o}),
    .b({_al_u863_o,\t/a/ID_rs1$0$_placeOpt_9 }),
    .c({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u867_o,\t/a/regfile/regfile$12$ [15]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [15]}),
    .mi({open_n22271,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u868_o,_al_u865_o}),
    .q({open_n22286,\t/a/regfile/regfile$12$ [15]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u878|t/a/regfile/reg0_b911  (
    .a({_al_u873_o,_al_u874_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .c({_al_u877_o,\t/a/ID_rs1$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u875_o,\t/a/regfile/regfile$28$ [15]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [15]}),
    .mi({open_n22288,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u878_o,_al_u875_o}),
    .q({open_n22303,\t/a/regfile/regfile$28$ [15]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u884 (
    .a({_al_u880_o,_al_u880_o}),
    .b({_al_u881_o,_al_u881_o}),
    .c({_al_u882_o,_al_u882_o}),
    .d({_al_u883_o,_al_u883_o}),
    .mi({open_n22316,\t/a/ID_rs1$2$_placeOpt_5 }),
    .fx({open_n22321,_al_u884_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u889|t/a/regfile/reg0_b398  (
    .a({_al_u884_o,_al_u885_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .c({_al_u888_o,\t/a/ID_rs1$1$_placeOpt_11 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u886_o,\t/a/regfile/regfile$12$ [14]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [14]}),
    .mi({open_n22325,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u889_o,_al_u886_o}),
    .q({open_n22340,\t/a/regfile/regfile$12$ [14]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u894 (
    .a({_al_u890_o,_al_u890_o}),
    .b({_al_u891_o,_al_u891_o}),
    .c({_al_u892_o,_al_u892_o}),
    .d({_al_u893_o,_al_u893_o}),
    .mi({open_n22353,\t/a/ID_rs1$2$_placeOpt_2 }),
    .fx({open_n22358,_al_u894_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u899|t/a/regfile/reg0_b910  (
    .a({_al_u894_o,_al_u895_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .c({_al_u898_o,\t/a/ID_rs1$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u896_o,\t/a/regfile/regfile$28$ [14]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [14]}),
    .mi({open_n22362,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u899_o,_al_u896_o}),
    .q({open_n22377,\t/a/regfile/regfile$28$ [14]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1000100010001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u910|t/a/regfile/reg0_b653  (
    .a({_al_u905_o,_al_u906_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .c({_al_u909_o,\t/a/ID_rs1$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u907_o,\t/a/regfile/regfile$20$ [13]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [13]}),
    .mi({open_n22379,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u910_o,_al_u907_o}),
    .q({open_n22394,\t/a/regfile/regfile$20$ [13]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110001011100),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u920|t/a/regfile/reg0_b397  (
    .a({_al_u917_o,_al_u916_o}),
    .b({_al_u915_o,\t/a/ID_rs1$0$_placeOpt_21 }),
    .c({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$1$_placeOpt_21 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u919_o,\t/a/regfile/regfile$12$ [13]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [13]}),
    .mi({open_n22396,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u920_o,_al_u917_o}),
    .q({open_n22411,\t/a/regfile/regfile$12$ [13]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u926 (
    .a({_al_u922_o,_al_u922_o}),
    .b({_al_u923_o,_al_u923_o}),
    .c({_al_u924_o,_al_u924_o}),
    .d({_al_u925_o,_al_u925_o}),
    .mi({open_n22424,\t/a/ID_rs1$2$_placeOpt_3 }),
    .fx({open_n22429,_al_u926_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u931|t/a/regfile/reg0_b396  (
    .a({_al_u926_o,_al_u927_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_1 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .c({_al_u930_o,\t/a/ID_rs1$1$_placeOpt_17 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u928_o,\t/a/regfile/regfile$12$ [12]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [12]}),
    .mi({open_n22433,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u931_o,_al_u928_o}),
    .q({open_n22448,\t/a/regfile/regfile$12$ [12]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u936 (
    .a({_al_u932_o,_al_u932_o}),
    .b({_al_u933_o,_al_u933_o}),
    .c({_al_u934_o,_al_u934_o}),
    .d({_al_u935_o,_al_u935_o}),
    .mi({open_n22461,\t/a/ID_rs1$2$_placeOpt_7 }),
    .fx({open_n22466,_al_u936_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(B*~((~D*~A))*~(C)+B*(~D*~A)*~(C)+~(B)*(~D*~A)*C+B*(~D*~A)*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000110001011100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u941|t/a/regfile/reg0_b908  (
    .a({_al_u938_o,_al_u937_o}),
    .b({_al_u936_o,\t/a/ID_rs1$0$_placeOpt_14 }),
    .c({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u940_o,\t/a/regfile/regfile$28$ [12]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [12]}),
    .mi({open_n22470,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u941_o,_al_u938_o}),
    .q({open_n22485,\t/a/regfile/regfile$28$ [12]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1000100010001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u952|t/a/regfile/reg0_b651  (
    .a({_al_u947_o,_al_u948_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .c({_al_u951_o,\t/a/ID_rs1$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u949_o,\t/a/regfile/regfile$20$ [11]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [11]}),
    .mi({open_n22487,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u952_o,_al_u949_o}),
    .q({open_n22502,\t/a/regfile/regfile$20$ [11]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u962|t/a/regfile/reg0_b395  (
    .a({_al_u957_o,_al_u958_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_21 }),
    .c({_al_u961_o,\t/a/ID_rs1$1$_placeOpt_21 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u959_o,\t/a/regfile/regfile$12$ [11]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [11]}),
    .mi({open_n22504,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u962_o,_al_u959_o}),
    .q({open_n22519,\t/a/regfile/regfile$12$ [11]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u968 (
    .a({_al_u964_o,_al_u964_o}),
    .b({_al_u965_o,_al_u965_o}),
    .c({_al_u966_o,_al_u966_o}),
    .d({_al_u967_o,_al_u967_o}),
    .mi({open_n22532,\t/a/ID_rs1$2$_placeOpt_7 }),
    .fx({open_n22537,_al_u968_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001000101110),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u973|t/a/regfile/reg0_b394  (
    .a({_al_u968_o,_al_u969_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .c({_al_u972_o,\t/a/ID_rs1$1$_placeOpt_11 }),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u970_o,\t/a/regfile/regfile$12$ [10]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [10]}),
    .mi({open_n22541,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u973_o,_al_u970_o}),
    .q({open_n22556,\t/a/regfile/regfile$12$ [10]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u978 (
    .a({_al_u974_o,_al_u974_o}),
    .b({_al_u975_o,_al_u975_o}),
    .c({_al_u976_o,_al_u976_o}),
    .d({_al_u977_o,_al_u977_o}),
    .mi({open_n22569,\t/a/ID_rs1$2$_placeOpt_7 }),
    .fx({open_n22574,_al_u978_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~D))*~(B)+A*(~C*~D)*~(B)+~(A)*(~C*~D)*B+A*(~C*~D)*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0010001000101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u983|t/a/regfile/reg0_b906  (
    .a({_al_u978_o,_al_u979_o}),
    .b({\t/a/ID_rs1$3$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .c({_al_u982_o,\t/a/ID_rs1$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u980_o,\t/a/regfile/regfile$28$ [10]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [10]}),
    .mi({open_n22578,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u983_o,_al_u980_o}),
    .q({open_n22593,\t/a/regfile/regfile$28$ [10]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*~C*~B*A)"),
    //.LUTF1("~D*~B*~A*~C+D*~B*~A*~C+~D*~B*A*~C+D*~B*A*~C+~D*~B*~A*C+~D*~B*A*C"),
    //.LUTG0("(~1*D*~C*~B*A)"),
    //.LUTG1("D*~B*~A*~C+D*~B*A*~C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u985|t/a/regfile/reg0_b128  (
    .a({open_n22594,_al_u254_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_10 ,\t/a/WB_rd [0]}),
    .c({\t/a/regfile/regfile$5$ [0],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$4$ [0],\t/a/WB_rd [3]}),
    .mi({open_n22596,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u985_o,\t/a/regfile/mux39_b128_sel_is_3_o }),
    .q({open_n22611,\t/a/regfile/regfile$4$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*C*~B*A)"),
    //.LUTF1("~A*C*~B*~D+A*C*~B*~D+~A*C*B*~D+A*C*B*~D+A*C*~B*D+A*C*B*D"),
    //.LUTG0("(~1*D*C*~B*A)"),
    //.LUTG1("~A*C*~B*~D+~A*C*B*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b1010000011110000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u986|t/a/regfile/reg0_b192  (
    .a({\t/a/ID_rs1$0$_placeOpt_16 ,_al_u254_o}),
    .b({open_n22612,\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$6$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$7$ [0],\t/a/WB_rd [3]}),
    .mi({open_n22614,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u986_o,\t/a/regfile/mux39_b192_sel_is_3_o }),
    .q({open_n22629,\t/a/regfile/regfile$6$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~A)*~((~B*~C))*~(0)+(~D*~A)*(~B*~C)*~(0)+~((~D*~A))*(~B*~C)*0+(~D*~A)*(~B*~C)*0)"),
    //.LUTF1("~A*~C*~D*~B+A*~C*~D*~B+A*~C*D*~B+~A*~C*~D*B+A*~C*~D*B+A*~C*D*B"),
    //.LUTG0("~((~D*~A)*~((~B*~C))*~(1)+(~D*~A)*(~B*~C)*~(1)+~((~D*~A))*(~B*~C)*1+(~D*~A)*(~B*~C)*1)"),
    //.LUTG1("~A*~C*~D*~B+~A*~C*~D*B"),
    .INIT_LUTF0(16'b1111111110101010),
    .INIT_LUTF1(16'b0000101000001111),
    .INIT_LUTG0(16'b1111110011111100),
    .INIT_LUTG1(16'b0000000000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u987|_al_u989  (
    .a({\t/a/ID_rs1$0$_placeOpt_16 ,_al_u987_o}),
    .b({open_n22630,_al_u986_o}),
    .c({\t/a/ID_rs1$1$_placeOpt_16 ,_al_u985_o}),
    .d({\t/a/regfile/regfile$0$ [0],_al_u988_o}),
    .e({\t/a/regfile/regfile$1$ [0],\t/a/ID_rs1$2$_placeOpt_6 }),
    .f({_al_u987_o,_al_u989_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u988|t/a/regfile/reg0_b96  (
    .a({\t/a/regfile/regfile$2$ [0],_al_u2614_o}),
    .b({\t/a/regfile/regfile$3$ [0],_al_u2616_o}),
    .c({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/MEM_aludat [0]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/reg_writedat [0]}),
    .mi({open_n22663,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u988_o,_al_u2760_o}),
    .q({open_n22667,\t/a/regfile/regfile$3$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u990|_al_u1706  (
    .a({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/ID_rs1$2$_placeOpt_6 ,\t/a/ID_rs2$2$_placeOpt_7 }),
    .d({\t/a/regfile/regfile$14$ [0],\t/a/regfile/regfile$14$ [0]}),
    .e({\t/a/regfile/regfile$15$ [0],\t/a/regfile/regfile$15$ [0]}),
    .f({_al_u990_o,_al_u1706_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*~B*A)"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(1*D*~C*~B*A)"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u991|t/a/regfile/reg0_b384  (
    .a({_al_u990_o,_al_u254_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/WB_rd [0]}),
    .c({\t/a/regfile/regfile$12$ [0],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$13$ [0],\t/a/WB_rd [3]}),
    .mi({open_n22691,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u991_o,\t/a/regfile/mux39_b384_sel_is_3_o }),
    .q({open_n22706,\t/a/regfile/regfile$12$ [0]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUT1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUT0(16'b0000011100000011),
    .INIT_LUT1(16'b0000111100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u992 (
    .a({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/ID_rs1$0$_placeOpt_16 }),
    .b({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/ID_rs1$1$_placeOpt_16 }),
    .c({\t/a/ID_rs1$2$_placeOpt_6 ,\t/a/ID_rs1$2$_placeOpt_6 }),
    .d({\t/a/regfile/regfile$10$ [0],\t/a/regfile/regfile$10$ [0]}),
    .mi({open_n22719,\t/a/regfile/regfile$11$ [0]}),
    .fx({open_n22724,_al_u992_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~D*~B))*~(C)+A*(~D*~B)*~(C)+~(A)*(~D*~B)*C+A*(~D*~B)*C))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~D*~B))*~(C)+A*(~D*~B)*~(C)+~(A)*(~D*~B)*C+A*(~D*~B)*C))"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000101000111010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u994|_al_u993  (
    .a({_al_u989_o,_al_u992_o}),
    .b({_al_u991_o,\t/a/ID_rs1$0$_placeOpt_16 }),
    .c({\t/a/ID_rs1 [3],\t/a/ID_rs1$1$_placeOpt_16 }),
    .d({_al_u993_o,\t/a/regfile/regfile$8$ [0]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$9$ [0]}),
    .f({_al_u994_o,_al_u993_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*~C*~B*A)"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D+~A*~C*B*~D+A*~C*B*~D+A*~C*~B*D+A*~C*B*D"),
    //.LUTG0("(~1*D*~C*~B*A)"),
    //.LUTG1("~A*~C*~B*~D+~A*~C*B*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000101000001111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u995|t/a/regfile/reg0_b640  (
    .a({\t/a/ID_rs1$0$_placeOpt_10 ,_al_u256_o}),
    .b({open_n22749,\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs1$1$_placeOpt_10 ,\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$20$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$21$ [0],\t/a/WB_rd [3]}),
    .mi({open_n22751,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u995_o,\t/a/regfile/mux39_b640_sel_is_3_o }),
    .q({open_n22766,\t/a/regfile/regfile$20$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~A*~B))*~(0)+(~D*~C)*(~A*~B)*~(0)+~((~D*~C))*(~A*~B)*0+(~D*~C)*(~A*~B)*0)"),
    //.LUTF1("~A*C*~B*~D+A*C*~B*~D+~A*C*B*~D+A*C*B*~D+~A*C*~B*D+~A*C*B*D"),
    //.LUTG0("~((~D*~C)*~((~A*~B))*~(1)+(~D*~C)*(~A*~B)*~(1)+~((~D*~C))*(~A*~B)*1+(~D*~C)*(~A*~B)*1)"),
    //.LUTG1("A*C*~B*~D+A*C*B*~D"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0101000011110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u996|_al_u999  (
    .a({\t/a/ID_rs1$0$_placeOpt_10 ,_al_u996_o}),
    .b({open_n22767,_al_u995_o}),
    .c({\t/a/ID_rs1$1$_placeOpt_10 ,_al_u997_o}),
    .d({\t/a/regfile/regfile$23$ [0],_al_u998_o}),
    .e({\t/a/regfile/regfile$22$ [0],\t/a/ID_rs1$2$_placeOpt_4 }),
    .f({_al_u996_o,_al_u999_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~D*~B+A*~C*~D*~B+A*~C*D*~B+~A*~C*~D*B+A*~C*~D*B+A*~C*D*B"),
    //.LUTF1("~C*~B*~D*~A+C*~B*~D*~A+C*~B*D*~A+~C*~B*~D*A+C*~B*~D*A+C*~B*D*A"),
    //.LUTG0("~A*~C*~D*~B+~A*~C*~D*B"),
    //.LUTG1("~C*~B*~D*~A+~C*~B*~D*A"),
    .INIT_LUTF0(16'b0000101000001111),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0000000000000101),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u997|_al_u1713  (
    .a({open_n22790,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/ID_rs1$1$_placeOpt_10 ,open_n22791}),
    .c({\t/a/ID_rs1$0$_placeOpt_10 ,\t/a/ID_rs2$1$_placeOpt_12 }),
    .d({\t/a/regfile/regfile$16$ [0],\t/a/regfile/regfile$16$ [0]}),
    .e({\t/a/regfile/regfile$17$ [0],\t/a/regfile/regfile$17$ [0]}),
    .f({_al_u997_o,_al_u1713_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"))
    \_al_u998|_al_u1714  (
    .a({\t/a/ID_rs1$0$_placeOpt_10 ,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/ID_rs1$1$_placeOpt_10 ,\t/a/ID_rs2$1$_placeOpt_12 }),
    .c({\t/a/regfile/regfile$18$ [0],\t/a/regfile/regfile$18$ [0]}),
    .d({\t/a/regfile/regfile$19$ [0],\t/a/regfile/regfile$19$ [0]}),
    .f({_al_u998_o,_al_u1714_o}));
  // address_offset=0;data_offset=0;depth=64;width=9;num_section=1;width_per_section=9;section_size=97;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    //.RID("0x0004"),
    //.WID("0x0004"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    auto_chipwatcher_0_logicbram_64x97_sub_000000_000 (
    .addra({4'b0000,status_5,status_4,status_3,status_2,status_1,status_0,3'b111}),
    .cea(wt_ce),
    .ceb(wt_ce),
    .clka(clock_pad),
    .dia({addr[17:10],addr[0]}),
    .wea(wt_ce),
    .web(wt_ce));
  // address_offset=0;data_offset=9;depth=64;width=9;num_section=1;width_per_section=9;section_size=97;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    //.RID("0x0005"),
    //.WID("0x0005"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    auto_chipwatcher_0_logicbram_64x97_sub_000000_009 (
    .addra({4'b0000,status_5,status_4,status_3,status_2,status_1,status_0,3'b111}),
    .cea(wt_ce),
    .ceb(wt_ce),
    .clka(clock_pad),
    .dia({addr[25:20],addr[1],addr[19:18]}),
    .wea(wt_ce),
    .web(wt_ce));
  // address_offset=0;data_offset=18;depth=64;width=9;num_section=1;width_per_section=9;section_size=97;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    //.RID("0x0006"),
    //.WID("0x0006"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    auto_chipwatcher_0_logicbram_64x97_sub_000000_018 (
    .addra({4'b0000,status_5,status_4,status_3,status_2,status_1,status_0,3'b111}),
    .cea(wt_ce),
    .ceb(wt_ce),
    .clka(clock_pad),
    .dia({addr[4:3],addr[31:30],addr[2],addr[29:26]}),
    .wea(wt_ce),
    .web(wt_ce));
  // address_offset=0;data_offset=27;depth=64;width=9;num_section=1;width_per_section=9;section_size=97;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    //.RID("0x0007"),
    //.WID("0x0007"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    auto_chipwatcher_0_logicbram_64x97_sub_000000_027 (
    .addra({4'b0000,status_5,status_4,status_3,status_2,status_1,status_0,3'b111}),
    .cea(wt_ce),
    .ceb(wt_ce),
    .clka(clock_pad),
    .dia({i_data[12:10],i_data[0],addr[9:5]}),
    .wea(wt_ce),
    .web(wt_ce));
  // address_offset=0;data_offset=36;depth=64;width=9;num_section=1;width_per_section=9;section_size=97;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    //.RID("0x0008"),
    //.WID("0x0008"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    auto_chipwatcher_0_logicbram_64x97_sub_000000_036 (
    .addra({4'b0000,status_5,status_4,status_3,status_2,status_1,status_0,3'b111}),
    .cea(wt_ce),
    .ceb(wt_ce),
    .clka(clock_pad),
    .dia({i_data[20],i_data[1],i_data[19:13]}),
    .wea(wt_ce),
    .web(wt_ce));
  // address_offset=0;data_offset=45;depth=64;width=9;num_section=1;width_per_section=9;section_size=97;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    //.RID("0x0009"),
    //.WID("0x0009"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    auto_chipwatcher_0_logicbram_64x97_sub_000000_045 (
    .addra({4'b0000,status_5,status_4,status_3,status_2,status_1,status_0,3'b111}),
    .cea(wt_ce),
    .ceb(wt_ce),
    .clka(clock_pad),
    .dia(i_data[29:21]),
    .wea(wt_ce),
    .web(wt_ce));
  // address_offset=0;data_offset=54;depth=64;width=9;num_section=1;width_per_section=9;section_size=97;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    //.RID("0x000A"),
    //.WID("0x000A"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    auto_chipwatcher_0_logicbram_64x97_sub_000000_054 (
    .addra({4'b0000,status_5,status_4,status_3,status_2,status_1,status_0,3'b111}),
    .cea(wt_ce),
    .ceb(wt_ce),
    .clka(clock_pad),
    .dia({i_data[8:3],i_data[31:30],i_data[2]}),
    .wea(wt_ce),
    .web(wt_ce));
  // address_offset=0;data_offset=63;depth=64;width=9;num_section=1;width_per_section=9;section_size=97;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    //.RID("0x000B"),
    //.WID("0x000B"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    auto_chipwatcher_0_logicbram_64x97_sub_000000_063 (
    .addra({4'b0000,status_5,status_4,status_3,status_2,status_1,status_0,3'b111}),
    .cea(wt_ce),
    .ceb(wt_ce),
    .clka(clock_pad),
    .dia({o_data[16:10],o_data[0],i_data[9]}),
    .wea(wt_ce),
    .web(wt_ce));
  // address_offset=0;data_offset=72;depth=64;width=9;num_section=1;width_per_section=9;section_size=97;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    //.RID("0x000C"),
    //.WID("0x000C"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    auto_chipwatcher_0_logicbram_64x97_sub_000000_072 (
    .addra({4'b0000,status_5,status_4,status_3,status_2,status_1,status_0,3'b111}),
    .cea(wt_ce),
    .ceb(wt_ce),
    .clka(clock_pad),
    .dia({o_data[24:20],o_data[1],o_data[19:17]}),
    .wea(wt_ce),
    .web(wt_ce));
  // address_offset=0;data_offset=81;depth=64;width=9;num_section=1;width_per_section=9;section_size=97;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    //.RID("0x000D"),
    //.WID("0x000D"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    auto_chipwatcher_0_logicbram_64x97_sub_000000_081 (
    .addra({4'b0000,status_5,status_4,status_3,status_2,status_1,status_0,3'b111}),
    .cea(wt_ce),
    .ceb(wt_ce),
    .clka(clock_pad),
    .dia({o_data[3],o_data[31:30],o_data[2],o_data[29:25]}),
    .wea(wt_ce),
    .web(wt_ce));
  // address_offset=0;data_offset=90;depth=64;width=7;num_section=1;width_per_section=7;section_size=97;working_depth=1024;working_width=9;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.FORCE_KEEP("ON"),
    //.RID("0x000E"),
    //.WID("0x000E"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("SP8K"),
    .OCEAMUX("1"),
    .OCEBMUX("1"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    auto_chipwatcher_0_logicbram_64x97_sub_000000_090 (
    .addra({4'b0000,status_5,status_4,status_3,status_2,status_1,status_0,3'b111}),
    .cea(wt_ce),
    .ceb(wt_ce),
    .clka(clock_pad),
    .dia({open_n23364,open_n23365,rst_pad,o_data[9:4]}),
    .wea(wt_ce),
    .web(wt_ce));
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(1)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*1*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111011011100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b0  (
    .a({_al_u3035_o,_al_u3034_o}),
    .b({_al_u3034_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [0],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [0]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [1],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [1]}),
    .mi({open_n23408,status_0}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23414,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [0]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(1)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*1*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111010111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b1  (
    .a({_al_u3034_o,_al_u3034_o}),
    .b({_al_u3035_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [1],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [1]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [2],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [2]}),
    .mi({open_n23426,status_1}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23432,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [1]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*~(1)*~(A)+(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*1*~(A)+~((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))*1*A+(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*1*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111101111101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b10  (
    .a({_al_u3034_o,_al_u3034_o}),
    .b({_al_u3035_o,_al_u3035_o}),
    .c(\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [11:10]),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [10],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [11]}),
    .mi({open_n23444,status_10}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23450,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [10]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(1)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*1*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111010111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b11  (
    .a({_al_u3034_o,_al_u3034_o}),
    .b({_al_u3035_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [11],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [11]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [12],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [12]}),
    .mi({open_n23462,status_11}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23468,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [11]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(1)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*1*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111010111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b12  (
    .a({_al_u3034_o,_al_u3034_o}),
    .b({_al_u3035_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [12],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [12]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [13],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [13]}),
    .mi({open_n23480,status_12}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23486,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [12]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*~(1)*~(A)+(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*1*~(A)+~((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))*1*A+(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*1*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111101111101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b13  (
    .a({_al_u3034_o,_al_u3034_o}),
    .b({_al_u3035_o,_al_u3035_o}),
    .c(\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [14:13]),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [13],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [14]}),
    .mi({open_n23498,status_13}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23504,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [13]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(1)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*1*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111010111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b14  (
    .a({_al_u3034_o,_al_u3034_o}),
    .b({_al_u3035_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [14],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [14]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [15],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [15]}),
    .mi({open_n23516,status_14}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23522,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [14]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(1)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*1*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111011011100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b15  (
    .a({_al_u3035_o,_al_u3034_o}),
    .b({_al_u3034_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [15],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [15]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [16],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [16]}),
    .mi({open_n23534,status_15}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23540,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [15]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(1)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*1*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111011011100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b16  (
    .a({_al_u3035_o,_al_u3034_o}),
    .b({_al_u3034_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [16],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [16]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [17],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [17]}),
    .mi({open_n23552,status_16}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23558,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [16]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(1)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*1*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111010111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b2  (
    .a({_al_u3034_o,_al_u3034_o}),
    .b({_al_u3035_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [2],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [2]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [3],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [3]}),
    .mi({open_n23570,status_2}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23576,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [2]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(1)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*1*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111011011100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b3  (
    .a({_al_u3035_o,_al_u3034_o}),
    .b({_al_u3034_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [3],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [3]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [4],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [4]}),
    .mi({open_n23588,status_3}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23594,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [3]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(1)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*1*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111010111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b4  (
    .a({_al_u3034_o,_al_u3034_o}),
    .b({_al_u3035_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [4],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [4]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [5],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [5]}),
    .mi({open_n23606,status_4}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23612,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [4]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(1)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*1*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111010111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b5  (
    .a({_al_u3034_o,_al_u3034_o}),
    .b({_al_u3035_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [5],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [5]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [6],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [6]}),
    .mi({open_n23624,status_5}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23630,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [5]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(1)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*1*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111011011100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b6  (
    .a({_al_u3035_o,_al_u3034_o}),
    .b({_al_u3034_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [6],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [6]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [7],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [7]}),
    .mi({open_n23642,status_6}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23648,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [6]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(1)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*1*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*1*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111010111010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b7  (
    .a({_al_u3034_o,_al_u3034_o}),
    .b({_al_u3035_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [7],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [7]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [8],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [8]}),
    .mi({open_n23660,status_7}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23666,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [7]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*~(0)*~(A)+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*~(A)+~((C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))*0*A+(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)*0*A)"),
    //.LUT1("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(1)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*1*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*1*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111111011011100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b8  (
    .a({_al_u3035_o,_al_u3034_o}),
    .b({_al_u3034_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [8],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [8]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [9],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [9]}),
    .mi({open_n23678,status_8}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23684,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [8]}));  // D:/td/td/cw\register.v(31)
  EG_PHY_MSLICE #(
    //.LUT0("((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*~(0)*~(A)+(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*0*~(A)+~((D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))*0*A+(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)*0*A)"),
    //.LUT1("((D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*~(1)*~(B)+(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*1*~(B)+~((D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))*1*B+(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)*1*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b1111110111101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg0_b9  (
    .a({_al_u3035_o,_al_u3034_o}),
    .b({_al_u3034_o,_al_u3035_o}),
    .c({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [10],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [10]}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [9],\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [9]}),
    .mi({open_n23696,status_9}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .q({open_n23702,\cfg_int/wrapper_cfg_inst/reg_inst/sshift_r2 [9]}));  // D:/td/td/cw\register.v(31)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b101|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b100  (
    .a({control_100,control_100}),
    .b({control_101,control_101}),
    .c({control_102,control_102}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [101:100]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3365_o,_al_u3366_o}),
    .q({control_101,control_100}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b102|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b33  (
    .a({_al_u3364_o,_al_u3308_o}),
    .b({_al_u3365_o,_al_u3309_o}),
    .c({control_102,_al_u3310_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3366_o,control_33}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [102],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [33]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3367_o,_al_u3311_o}),
    .q({control_102,control_33}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b104|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b103  (
    .a({control_103,control_103}),
    .b({control_104,control_104}),
    .c({control_105,control_105}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [104:103]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3348_o,_al_u3349_o}),
    .q({control_104,control_103}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b105|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b303  (
    .a({_al_u3347_o,_al_u3382_o}),
    .b({_al_u3348_o,_al_u3383_o}),
    .c({_al_u3349_o,_al_u3384_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_105,control_303}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [105],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [303]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3350_o,_al_u3385_o}),
    .q({control_105,control_303}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b107|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b106  (
    .a({control_106,control_106}),
    .b({control_107,control_107}),
    .c({control_108,control_108}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [107:106]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3353_o,_al_u3354_o}),
    .q({control_107,control_106}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b108|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b30  (
    .a({_al_u3352_o,_al_u3454_o}),
    .b({_al_u3353_o,_al_u3455_o}),
    .c({control_108,_al_u3456_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3354_o,control_30}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [108],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [30]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3355_o,_al_u3457_o}),
    .q({control_108,control_30}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b10|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b9  (
    .ce(jupdate),
    .clk(jtck),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [10:9]),
    .sr(\cfg_int/wrapper_cfg_inst/rst ),
    .q({control_10,control_9}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b110|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b109  (
    .a({control_109,control_109}),
    .b({control_110,control_110}),
    .c({control_111,control_111}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [110:109]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3374_o,_al_u3375_o}),
    .q({control_110,control_109}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b111|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b291  (
    .a({_al_u3373_o,_al_u3394_o}),
    .b({_al_u3374_o,_al_u3395_o}),
    .c({_al_u3375_o,_al_u3396_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_111,control_291}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [111],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [291]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3376_o,_al_u3397_o}),
    .q({control_111,control_291}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b113|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b112  (
    .a({control_112,control_112}),
    .b({control_113,control_113}),
    .c({control_114,control_114}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [113:112]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .f({_al_u3224_o,_al_u3225_o}),
    .q({control_113,control_112}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b114|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b285  (
    .a({_al_u3223_o,_al_u3509_o}),
    .b({_al_u3224_o,_al_u3510_o}),
    .c({control_114,_al_u3511_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3225_o,control_285}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [114],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [285]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .f({_al_u3226_o,_al_u3512_o}),
    .q({control_114,control_285}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b116|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b115  (
    .a({control_115,control_115}),
    .b({control_116,control_116}),
    .c({control_117,control_117}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [116:115]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3207_o,_al_u3208_o}),
    .q({control_116,control_115}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b117|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b279  (
    .a({_al_u3206_o,_al_u3424_o}),
    .b({_al_u3207_o,_al_u3425_o}),
    .c({control_117,_al_u3426_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3208_o,control_279}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [117],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [279]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3209_o,_al_u3427_o}),
    .q({control_117,control_279}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b119|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b118  (
    .a({control_118,control_118}),
    .b({control_119,control_119}),
    .c({control_120,control_120}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [119:118]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3211_o,_al_u3212_o}),
    .q({control_119,control_118}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b11|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b21  (
    .ce(jupdate),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [11],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [21]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_1 ),
    .q({control_11,control_21}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b120|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b270  (
    .a({_al_u3210_o,_al_u3420_o}),
    .b({_al_u3211_o,_al_u3421_o}),
    .c({_al_u3212_o,_al_u3422_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_120,control_270}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [120],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [270]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3213_o,_al_u3423_o}),
    .q({control_120,control_270}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b122|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b121  (
    .a({control_121,control_121}),
    .b({control_122,control_122}),
    .c({control_123,control_123}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [122:121]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .f({_al_u3228_o,_al_u3229_o}),
    .q({control_122,control_121}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b123|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b267  (
    .a({_al_u3227_o,_al_u3501_o}),
    .b({_al_u3228_o,_al_u3502_o}),
    .c({control_123,_al_u3503_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3229_o,control_267}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [123],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [267]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .f({_al_u3230_o,_al_u3504_o}),
    .q({control_123,control_267}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b125|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b124  (
    .a({control_124,control_124}),
    .b({control_125,control_125}),
    .c({control_126,control_126}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [125:124]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3370_o,_al_u3371_o}),
    .q({control_125,control_124}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b126|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b261  (
    .a({_al_u3369_o,_al_u3287_o}),
    .b({_al_u3370_o,_al_u3288_o}),
    .c({_al_u3371_o,_al_u3289_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_126,control_261}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [126],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [261]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3372_o,_al_u3290_o}),
    .q({control_126,control_261}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b128|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b127  (
    .a({control_127,control_127}),
    .b({control_128,control_128}),
    .c({control_129,control_129}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [128:127]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3254_o,_al_u3255_o}),
    .q({control_128,control_127}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b129|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b258  (
    .a({_al_u3253_o,_al_u3496_o}),
    .b({_al_u3254_o,_al_u3497_o}),
    .c({control_129,_al_u3498_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3255_o,control_258}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [129],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [258]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3256_o,_al_u3499_o}),
    .q({control_129,control_258}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b12|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b20  (
    .ce(jupdate),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [12],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [20]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_15 ),
    .q({control_12,control_20}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b131|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b130  (
    .a({control_130,control_130}),
    .b({control_131,control_131}),
    .c({control_132,control_132}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [131:130]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3233_o,_al_u3234_o}),
    .q({control_131,control_130}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b132|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b252  (
    .a({_al_u3232_o,_al_u3167_o}),
    .b({_al_u3233_o,_al_u3168_o}),
    .c({_al_u3234_o,_al_u3169_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_132,control_252}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [132],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [252]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3235_o,_al_u3170_o}),
    .q({control_132,control_252}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b134|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b133  (
    .a({control_133,control_133}),
    .b({control_134,control_134}),
    .c({control_135,control_135}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [134:133]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3216_o,_al_u3217_o}),
    .q({control_134,control_133}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b135|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b243  (
    .a({_al_u3215_o,_al_u3283_o}),
    .b({_al_u3216_o,_al_u3284_o}),
    .c({_al_u3217_o,_al_u3285_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_135,control_243}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [135],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [243]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3218_o,_al_u3286_o}),
    .q({control_135,control_243}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b137|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b136  (
    .a({control_136,control_136}),
    .b({control_137,control_137}),
    .c({control_138,control_138}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [137:136]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3340_o,_al_u3341_o}),
    .q({control_137,control_136}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b138|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b240  (
    .a({_al_u3339_o,_al_u3125_o}),
    .b({_al_u3340_o,_al_u3126_o}),
    .c({_al_u3341_o,_al_u3127_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_138,control_240}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [138],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [240]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3342_o,_al_u3128_o}),
    .q({control_138,control_240}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b13|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b19  (
    .ce(jupdate),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [13],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [19]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_15 ),
    .q({control_13,control_19}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b140|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b139  (
    .a({control_140,control_139}),
    .b({control_139,control_140}),
    .c({control_141,control_141}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [140:139]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3472_o,_al_u3473_o}),
    .q({control_140,control_139}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b141|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b24  (
    .a({_al_u3471_o,_al_u3180_o}),
    .b({_al_u3472_o,_al_u3181_o}),
    .c({control_141,_al_u3182_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3473_o,control_24}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [141],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [24]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3474_o,_al_u3183_o}),
    .q({control_141,control_24}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b143|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b142  (
    .a({control_142,control_142}),
    .b({control_143,control_143}),
    .c({control_144,control_144}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [143:142]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3476_o,_al_u3477_o}),
    .q({control_143,control_142}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b144|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b237  (
    .a({_al_u3475_o,_al_u3121_o}),
    .b({_al_u3476_o,_al_u3122_o}),
    .c({control_144,_al_u3123_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3477_o,control_237}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [144],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [237]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3478_o,_al_u3124_o}),
    .q({control_144,control_237}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b146|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b145  (
    .a({control_145,control_145}),
    .b({control_146,control_146}),
    .c({control_147,control_147}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [146:145]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3344_o,_al_u3345_o}),
    .q({control_146,control_145}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b147|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b234  (
    .a({_al_u3343_o,_al_u3399_o}),
    .b({_al_u3344_o,_al_u3400_o}),
    .c({control_147,_al_u3401_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3345_o,control_234}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [147],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [234]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3346_o,_al_u3402_o}),
    .q({control_147,control_234}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b149|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b148  (
    .a({control_148,control_148}),
    .b({control_149,control_149}),
    .c({control_150,control_150}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [149:148]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .f({_al_u3237_o,_al_u3238_o}),
    .q({control_149,control_148}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b14|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b18  (
    .ce(jupdate),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [14],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [18]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_1 ),
    .q({control_14,control_18}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b150|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b225  (
    .a({_al_u3236_o,_al_u3325_o}),
    .b({_al_u3237_o,_al_u3326_o}),
    .c({_al_u3238_o,_al_u3327_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_150,control_225}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [150],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [225]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .f({_al_u3239_o,_al_u3328_o}),
    .q({control_150,control_225}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b152|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b151  (
    .a({control_151,control_151}),
    .b({control_152,control_152}),
    .c({control_153,control_153}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [152:151]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3220_o,_al_u3221_o}),
    .q({control_152,control_151}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b153|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b207  (
    .a({_al_u3219_o,_al_u3274_o}),
    .b({_al_u3220_o,_al_u3275_o}),
    .c({control_153,_al_u3276_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3221_o,control_207}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [153],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [207]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3222_o,_al_u3277_o}),
    .q({control_153,control_207}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b155|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b154  (
    .a({control_154,control_154}),
    .b({control_155,control_155}),
    .c({control_156,control_156}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [155:154]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3318_o,_al_u3319_o}),
    .q({control_155,control_154}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b156|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b204  (
    .a({_al_u3317_o,_al_u3488_o}),
    .b({_al_u3318_o,_al_u3489_o}),
    .c({_al_u3319_o,_al_u3490_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_156,control_204}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [156],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [204]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .f({_al_u3320_o,_al_u3491_o}),
    .q({control_156,control_204}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b158|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b157  (
    .a({control_157,control_157}),
    .b({control_158,control_158}),
    .c({control_159,control_159}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [158:157]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_13 ),
    .f({_al_u3113_o,_al_u3114_o}),
    .q({control_158,control_157}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b159|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b201  (
    .a({_al_u3112_o,_al_u3159_o}),
    .b({_al_u3113_o,_al_u3160_o}),
    .c({_al_u3114_o,_al_u3161_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_159,control_201}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [159],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [201]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_13 ),
    .f({_al_u3115_o,_al_u3162_o}),
    .q({control_159,control_201}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b15|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b17  (
    .ce(jupdate),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [15],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [17]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_15 ),
    .q({control_15,control_17}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b161|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b160  (
    .a({control_160,control_160}),
    .b({control_161,control_161}),
    .c({control_162,control_162}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [161:160]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3194_o,_al_u3195_o}),
    .q({control_161,control_160}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b162|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b198  (
    .a({_al_u3193_o,_al_u3416_o}),
    .b({_al_u3194_o,_al_u3417_o}),
    .c({control_162,_al_u3418_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3195_o,control_198}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [162],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [198]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3196_o,_al_u3419_o}),
    .q({control_162,control_198}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b164|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b163  (
    .a({control_163,control_163}),
    .b({control_164,control_164}),
    .c({control_165,control_165}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [164:163]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3130_o,_al_u3131_o}),
    .q({control_164,control_163}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b165|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b195  (
    .a({_al_u3129_o,_al_u3150_o}),
    .b({_al_u3130_o,_al_u3151_o}),
    .c({_al_u3131_o,_al_u3152_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_165,control_195}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [165],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [195]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3132_o,_al_u3153_o}),
    .q({control_165,control_195}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b167|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b166  (
    .a({control_166,control_166}),
    .b({control_167,control_167}),
    .c({control_168,control_168}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [167:166]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3105_o,_al_u3106_o}),
    .q({control_167,control_166}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~C*~(1*~(~B*~(~D*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000001100000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b168|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b192  (
    .a({_al_u3104_o,_al_u3198_o}),
    .b({_al_u3105_o,_al_u3199_o}),
    .c({_al_u3106_o,_al_u3200_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_168,control_192}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [168],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [192]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3107_o,_al_u3201_o}),
    .q({control_168,control_192}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b170|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b169  (
    .a({control_169,control_169}),
    .b({control_170,control_170}),
    .c({control_171,control_171}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [170:169]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3434_o,_al_u3435_o}),
    .q({control_170,control_169}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b171|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b189  (
    .a({_al_u3433_o,_al_u3278_o}),
    .b({_al_u3434_o,_al_u3279_o}),
    .c({control_171,_al_u3280_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3435_o,control_189}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [171],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [189]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3436_o,_al_u3281_o}),
    .q({control_171,control_189}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b173|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b172  (
    .a({control_172,control_172}),
    .b({control_173,control_173}),
    .c({control_174,control_174}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [173:172]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3468_o,_al_u3469_o}),
    .q({control_173,control_172}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b174|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b186  (
    .a({_al_u3467_o,_al_u3146_o}),
    .b({_al_u3468_o,_al_u3147_o}),
    .c({control_174,_al_u3148_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3469_o,control_186}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [174],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [186]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3470_o,_al_u3149_o}),
    .q({control_174,control_186}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b176|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b175  (
    .a({control_175,control_175}),
    .b({control_176,control_176}),
    .c({control_177,control_177}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [176:175]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3336_o,_al_u3337_o}),
    .q({control_176,control_175}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~(~B*~(~D*~A))))"),
    //.LUTF1("(~D*~(0*~(~B*~(~C*~A))))"),
    //.LUTG0("(~C*~(1*~(~B*~(~D*~A))))"),
    //.LUTG1("(~D*~(1*~(~B*~(~C*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001111),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0000001100000010),
    .INIT_LUTG1(16'b0000000000110010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b177|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b183  (
    .a({_al_u3335_o,_al_u3261_o}),
    .b({_al_u3336_o,_al_u3262_o}),
    .c({control_177,_al_u3263_o}),
    .ce(jupdate),
    .clk(jtck),
    .d({_al_u3337_o,control_183}),
    .e({\trig_node/trigger_node_int_0/force_acq_fin ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [177],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [183]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3338_o,_al_u3264_o}),
    .q({control_177,control_183}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b179|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b178  (
    .a({control_178,control_178}),
    .b({control_179,control_179}),
    .c({\trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/ctl_last ,control_180}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_180,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [179:178]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3438_o,_al_u3439_o}),
    .q({control_179,control_178}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b182|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b181  (
    .a({control_182,control_181}),
    .b({control_181,control_182}),
    .c({control_183,control_183}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [182:181]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3262_o,_al_u3263_o}),
    .q({control_182,control_181}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b185|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b184  (
    .a({control_185,control_184}),
    .b({control_184,control_185}),
    .c({control_186,control_186}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [185:184]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3147_o,_al_u3148_o}),
    .q({control_185,control_184}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b188|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b187  (
    .a({control_188,control_187}),
    .b({control_187,control_188}),
    .c({control_189,control_189}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [188:187]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3279_o,_al_u3280_o}),
    .q({control_188,control_187}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b191|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b190  (
    .a({control_191,control_190}),
    .b({control_190,control_191}),
    .c({control_192,control_192}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [191:190]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3199_o,_al_u3200_o}),
    .q({control_191,control_190}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b194|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b193  (
    .a({control_193,control_193}),
    .b({control_194,control_194}),
    .c({control_195,control_195}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [194:193]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3151_o,_al_u3152_o}),
    .q({control_194,control_193}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b197|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b196  (
    .a({control_197,control_196}),
    .b({control_196,control_197}),
    .c({control_198,control_198}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [197:196]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3417_o,_al_u3418_o}),
    .q({control_197,control_196}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b1|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b16  (
    .ce(jupdate),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [1],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [16]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_15 ),
    .q({control_1,control_16}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b200|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b199  (
    .a({control_200,control_199}),
    .b({control_199,control_200}),
    .c({control_201,control_201}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [200:199]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_13 ),
    .f({_al_u3160_o,_al_u3161_o}),
    .q({control_200,control_199}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b203|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b202  (
    .a({control_203,control_202}),
    .b({control_202,control_203}),
    .c({control_204,control_204}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [203:202]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3489_o,_al_u3490_o}),
    .q({control_203,control_202}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b206|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b205  (
    .a({control_205,control_205}),
    .b({control_206,control_206}),
    .c({\trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/ctl_last ,control_207}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_207,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [206:205]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3275_o,_al_u3276_o}),
    .q({control_206,control_205}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b209|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b208  (
    .a({control_208,control_208}),
    .b({control_209,control_209}),
    .c({control_210,control_210}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [209:208]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3203_o,_al_u3204_o}),
    .q({control_209,control_208}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b212|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b211  (
    .a({control_211,control_211}),
    .b({control_212,control_212}),
    .c({\trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/ctl_last ,control_213}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_213,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [212:211]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .f({_al_u3241_o,_al_u3242_o}),
    .q({control_212,control_211}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b215|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b214  (
    .a({control_214,control_214}),
    .b({control_215,control_215}),
    .c({\trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/ctl_last ,control_216}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_216,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [215:214]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .f({_al_u3245_o,_al_u3246_o}),
    .q({control_215,control_214}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b218|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b217  (
    .a({control_218,control_217}),
    .b({control_217,control_218}),
    .c({control_219,control_219}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [218:217]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3357_o,_al_u3358_o}),
    .q({control_218,control_217}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b221|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b220  (
    .a({control_221,control_220}),
    .b({control_220,control_221}),
    .c({control_222,control_222}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [221:220]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3493_o,_al_u3494_o}),
    .q({control_221,control_220}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b224|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b223  (
    .a({control_223,control_223}),
    .b({control_224,control_224}),
    .c({\trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/ctl_last ,control_225}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_225,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [224:223]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .f({_al_u3326_o,_al_u3327_o}),
    .q({control_224,control_223}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b227|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b226  (
    .a({control_227,control_226}),
    .b({control_226,control_227}),
    .c({control_228,control_228}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [227:226]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3330_o,_al_u3331_o}),
    .q({control_227,control_226}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b230|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b229  (
    .a({control_229,control_229}),
    .b({control_230,control_230}),
    .c({\trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/ctl_last ,control_231}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_231,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$69$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [230:229]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .f({_al_u3250_o,_al_u3251_o}),
    .q({control_230,control_229}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b233|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b232  (
    .a({control_232,control_232}),
    .b({control_233,control_233}),
    .c({control_234,control_234}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [233:232]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3400_o,_al_u3401_o}),
    .q({control_233,control_232}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b236|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b235  (
    .a({control_235,control_235}),
    .b({control_236,control_236}),
    .c({control_237,control_237}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [236:235]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3122_o,_al_u3123_o}),
    .q({control_236,control_235}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b239|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b238  (
    .a({control_239,control_238}),
    .b({control_238,control_239}),
    .c({control_240,control_240}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [239:238]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3126_o,_al_u3127_o}),
    .q({control_239,control_238}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b23|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b22  (
    .a({control_22,control_22}),
    .b({control_23,control_23}),
    .c({control_24,control_24}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [23:22]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3181_o,_al_u3182_o}),
    .q({control_23,control_22}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b242|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b241  (
    .a({control_242,control_241}),
    .b({control_241,control_242}),
    .c({control_243,control_243}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [242:241]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3284_o,_al_u3285_o}),
    .q({control_242,control_241}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b245|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b244  (
    .a({control_244,control_244}),
    .b({control_245,control_245}),
    .c({control_246,control_246}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [245:244]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_13 ),
    .f({_al_u3143_o,_al_u3144_o}),
    .q({control_245,control_244}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b248|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b247  (
    .a({control_247,control_247}),
    .b({control_248,control_248}),
    .c({control_249,control_249}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [248:247]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3164_o,_al_u3165_o}),
    .q({control_248,control_247}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b251|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b250  (
    .a({control_250,control_250}),
    .b({control_251,control_251}),
    .c({control_252,control_252}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [251:250]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3168_o,_al_u3169_o}),
    .q({control_251,control_250}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b254|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b253  (
    .a({control_253,control_253}),
    .b({control_254,control_254}),
    .c({\trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/ctl_last ,control_255}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_255,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [254:253]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3480_o,_al_u3481_o}),
    .q({control_254,control_253}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b257|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b256  (
    .a({control_257,control_256}),
    .b({control_256,control_257}),
    .c({control_258,control_258}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [257:256]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3497_o,_al_u3498_o}),
    .q({control_257,control_256}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b260|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b259  (
    .a({control_259,control_259}),
    .b({control_260,control_260}),
    .c({control_261,control_261}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [260:259]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3288_o,_al_u3289_o}),
    .q({control_260,control_259}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b263|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b262  (
    .a({control_263,control_262}),
    .b({control_262,control_263}),
    .c({control_264,control_264}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [263:262]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .f({_al_u3271_o,_al_u3272_o}),
    .q({control_263,control_262}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b266|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b265  (
    .a({control_266,control_265}),
    .b({control_265,control_266}),
    .c({control_267,control_267}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [266:265]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .f({_al_u3502_o,_al_u3503_o}),
    .q({control_266,control_265}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b269|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b268  (
    .a({control_268,control_268}),
    .b({control_269,control_269}),
    .c({\trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/ctl_last ,control_270}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_270,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [269:268]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3421_o,_al_u3422_o}),
    .q({control_269,control_268}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b26|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b25  (
    .a({control_25,control_25}),
    .b({control_26,control_26}),
    .c({control_27,control_27}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [26:25]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3258_o,_al_u3259_o}),
    .q({control_26,control_25}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b272|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b271  (
    .a({control_271,control_271}),
    .b({control_272,control_272}),
    .c({control_273,control_273}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [272:271]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3485_o,_al_u3486_o}),
    .q({control_272,control_271}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b275|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b274  (
    .a({control_275,control_274}),
    .b({control_274,control_275}),
    .c({control_276,control_276}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [275:274]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3156_o,_al_u3157_o}),
    .q({control_275,control_274}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b278|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b277  (
    .a({control_278,control_277}),
    .b({control_277,control_278}),
    .c({control_279,control_279}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [278:277]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3425_o,_al_u3426_o}),
    .q({control_278,control_277}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b281|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b280  (
    .a({control_281,control_280}),
    .b({control_280,control_281}),
    .c({control_282,control_282}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [281:280]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3267_o,_al_u3268_o}),
    .q({control_281,control_280}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b284|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b283  (
    .a({control_284,control_283}),
    .b({control_283,control_284}),
    .c({control_285,control_285}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [284:283]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .f({_al_u3510_o,_al_u3511_o}),
    .q({control_284,control_283}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b287|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b286  (
    .a({control_287,control_286}),
    .b({control_286,control_287}),
    .c({control_288,control_288}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [287:286]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3506_o,_al_u3507_o}),
    .q({control_287,control_286}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b290|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b289  (
    .a({control_289,control_289}),
    .b({control_290,control_290}),
    .c({\trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/ctl_last ,control_291}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_291,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [290:289]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3395_o,_al_u3396_o}),
    .q({control_290,control_289}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b293|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b292  (
    .a({control_292,control_292}),
    .b({control_293,control_293}),
    .c({control_294,control_294}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [293:292]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3514_o,_al_u3515_o}),
    .q({control_293,control_292}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b296|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b295  (
    .a({control_295,control_295}),
    .b({control_296,control_296}),
    .c({control_297,control_297}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [296:295]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3408_o,_al_u3409_o}),
    .q({control_296,control_295}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b299|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b298  (
    .a({control_298,control_298}),
    .b({control_299,control_299}),
    .c({\trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/ctl_last ,control_300}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_300,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [299:298]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3412_o,_al_u3413_o}),
    .q({control_299,control_298}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b29|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b28  (
    .a({control_28,control_28}),
    .b({control_29,control_29}),
    .c({control_30,control_30}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [29:28]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3455_o,_al_u3456_o}),
    .q({control_29,control_28}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_MSLICE #(
    //.LUT0("(B*D)"),
    //.LUT1("(~D*A*~(B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110000000000),
    .INIT_LUT1(16'b0000000000101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b2|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b0  (
    .a({control_2,open_n25320}),
    .b({_al_u3518_o,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [0]}),
    .c({_al_u3334_o,open_n25321}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_3,\cfg_int/wrapper_cfg_inst/shift_0 }),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [2],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [0]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .f({_al_u3519_o,jtdo_0}),
    .q({control_2,control_0}));  // D:/td/td/cw\register.v(38)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b3  (
    .ce(jupdate),
    .clk(jtck),
    .mi({open_n25353,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [3]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({open_n25359,control_3}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b302|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b301  (
    .a({control_301,control_301}),
    .b({control_302,control_302}),
    .c({\trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/ctl_last ,control_303}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_303,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [302:301]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3383_o,_al_u3384_o}),
    .q({control_302,control_301}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b305|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b304  (
    .a({control_305,control_304}),
    .b({control_304,control_305}),
    .c({control_306,control_306}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [305:304]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3387_o,_al_u3388_o}),
    .q({control_305,control_304}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b308|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b307  (
    .a({control_307,control_307}),
    .b({control_308,control_308}),
    .c({\trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/ctl_last ,control_309}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_309,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [308:307]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3404_o,_al_u3405_o}),
    .q({control_308,control_307}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b311|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b310  (
    .a({control_310,control_310}),
    .b({control_311,control_311}),
    .c({\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last ,control_312}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_312,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [311:310]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3391_o,_al_u3392_o}),
    .q({control_311,control_310}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b32|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b31  (
    .a({control_31,control_31}),
    .b({control_32,control_32}),
    .c({control_33,control_33}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [32:31]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3309_o,_al_u3310_o}),
    .q({control_32,control_31}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b35|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b34  (
    .a({control_35,control_34}),
    .b({control_34,control_35}),
    .c({control_36,control_36}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [35:34]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3313_o,_al_u3314_o}),
    .q({control_35,control_34}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b38|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b37  (
    .a({control_37,control_37}),
    .b({control_38,control_38}),
    .c({control_39,control_39}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [38:37]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .f({_al_u3459_o,_al_u3460_o}),
    .q({control_38,control_37}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b41|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b40  (
    .a({control_40,control_40}),
    .b({control_41,control_41}),
    .c({\trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/ctl_last ,control_42}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_42,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }),
    .e({\trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [41:40]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .f({_al_u3446_o,_al_u3447_o}),
    .q({control_41,control_40}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b44|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b43  (
    .a({control_43,control_43}),
    .b({control_44,control_44}),
    .c({control_45,control_45}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [44:43]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3429_o,_al_u3430_o}),
    .q({control_44,control_43}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~A*~B*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~A*~B*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b47|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b46  (
    .a({control_47,control_46}),
    .b({control_46,control_47}),
    .c({control_48,control_48}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [47:46]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3185_o,_al_u3186_o}),
    .q({control_47,control_46}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b50|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b49  (
    .a({control_49,control_49}),
    .b({control_50,control_50}),
    .c({\trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/ctl_last ,control_51}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_51,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [50:49]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .f({_al_u3322_o,_al_u3323_o}),
    .q({control_50,control_49}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b53|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b52  (
    .a({control_52,control_52}),
    .b({control_53,control_53}),
    .c({control_54,control_54}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [53:52]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3117_o,_al_u3118_o}),
    .q({control_53,control_52}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b56|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b55  (
    .a({control_55,control_55}),
    .b({control_56,control_56}),
    .c({control_57,control_57}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [56:55]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3463_o,_al_u3464_o}),
    .q({control_56,control_55}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b59|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b58  (
    .a({control_58,control_58}),
    .b({control_59,control_59}),
    .c({control_60,control_60}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [59:58]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3134_o,_al_u3135_o}),
    .q({control_59,control_58}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b62|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b61  (
    .a({control_61,control_61}),
    .b({control_62,control_62}),
    .c({control_63,control_63}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [62:61]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3177_o,_al_u3178_o}),
    .q({control_62,control_61}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b65|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b64  (
    .a({control_64,control_64}),
    .b({control_65,control_65}),
    .c({control_66,control_66}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [65:64]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3305_o,_al_u3306_o}),
    .q({control_65,control_64}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b68|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b67  (
    .a({control_67,control_67}),
    .b({control_68,control_68}),
    .c({control_69,control_69}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [68:67]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3451_o,_al_u3452_o}),
    .q({control_68,control_67}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b71|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b70  (
    .a({control_70,control_70}),
    .b({control_71,control_71}),
    .c({control_72,control_72}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [71:70]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3190_o,_al_u3191_o}),
    .q({control_71,control_70}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b74|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b73  (
    .a({control_73,control_73}),
    .b({control_74,control_74}),
    .c({control_75,control_75}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [74:73]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3139_o,_al_u3140_o}),
    .q({control_74,control_73}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b77|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b76  (
    .a({control_76,control_76}),
    .b({control_77,control_77}),
    .c({control_78,control_78}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [77:76]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .f({_al_u3292_o,_al_u3293_o}),
    .q({control_77,control_76}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b80|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b79  (
    .a({control_79,control_79}),
    .b({control_80,control_80}),
    .c({control_81,control_81}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [80:79]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .f({_al_u3442_o,_al_u3443_o}),
    .q({control_80,control_79}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b83|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b82  (
    .a({control_82,control_82}),
    .b({control_83,control_83}),
    .c({control_84,control_84}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [83:82]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .f({_al_u3301_o,_al_u3302_o}),
    .q({control_83,control_82}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b86|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b85  (
    .a({control_85,control_85}),
    .b({control_86,control_86}),
    .c({control_87,control_87}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }),
    .e({\trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [86:85]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .f({_al_u3296_o,_al_u3297_o}),
    .q({control_86,control_85}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b89|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b88  (
    .a({control_88,control_88}),
    .b({control_89,control_89}),
    .c({control_90,control_90}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }),
    .e({\trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [89:88]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .f({_al_u3173_o,_al_u3174_o}),
    .q({control_89,control_88}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b92|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b91  (
    .a({control_91,control_91}),
    .b({control_92,control_92}),
    .c({control_93,control_93}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }),
    .e({\trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [92:91]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .f({_al_u3109_o,_al_u3110_o}),
    .q({control_92,control_91}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(C*D*~(0)+~(C)*~(D)*0+C*~(D)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(C*D*~(1)+~(C)*~(D)*1+C*~(D)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b95|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b94  (
    .a({control_94,control_94}),
    .b({control_95,control_95}),
    .c({control_96,control_96}),
    .ce(jupdate),
    .clk(jtck),
    .d({\trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [95:94]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3361_o,_al_u3362_o}),
    .q({control_95,control_94}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(38)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(~B*~A*(D*C*~(0)+~(D)*~(C)*0+D*~(C)*0))"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(~B*~A*(D*C*~(1)+~(D)*~(C)*1+D*~(C)*1))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg1_b98|cfg_int/wrapper_cfg_inst/reg_inst/reg1_b97  (
    .a({control_97,control_97}),
    .b({control_98,control_98}),
    .c({\trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/ctl_last ,control_99}),
    .ce(jupdate),
    .clk(jtck),
    .d({control_99,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }),
    .e({\trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 }),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [98:97]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .f({_al_u3378_o,_al_u3379_o}),
    .q({control_98,control_97}));  // D:/td/td/cw\register.v(38)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b100|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b101  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [101],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [102]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [100],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [101]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b102|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b103  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [103],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [104]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [102],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [103]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b104|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b105  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [105],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [106]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [104],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [105]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b106|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b107  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [107],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [108]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [106],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [107]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b108|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b109  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [109],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [110]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [108],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [109]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b10|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b11  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [11],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [12]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_1 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [10],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [11]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b110|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b111  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [111],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [112]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [110],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [111]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b112|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b113  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [113],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [114]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [112],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [113]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b114|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b115  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [115],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [116]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [114],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [115]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b116|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b117  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [117],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [118]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [116],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [117]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b118|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b119  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [119],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [120]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [118],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [119]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b120|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b121  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [121],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [122]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [120],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [121]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b122|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b123  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [123],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [124]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [122],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [123]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b124|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b125  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [125],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [126]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [124],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [125]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b126|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b127  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [127],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [128]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [126],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [127]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b128|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b129  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [129],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [130]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [128],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [129]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b12|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b13  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [13],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [14]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_1 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [12],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [13]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b130|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b131  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [131],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [132]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [130],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [131]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b132|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b133  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [133],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [134]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [132],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [133]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b134|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b135  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [135],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [136]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [134],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [135]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b136|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b137  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [137],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [138]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [136],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [137]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b138|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b139  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [139],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [140]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [138],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [139]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b140|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b141  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [141],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [142]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [140],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [141]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b142|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b143  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [143],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [144]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_13 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [142],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [143]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b144|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b145  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [145],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [146]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [144],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [145]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b146|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b147  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [147],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [148]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [146],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [147]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b148|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b149  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [149],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [150]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [148],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [149]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b14|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b15  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [15],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [16]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_15 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [14],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [15]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b150|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b151  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [151],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [152]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [150],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [151]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b152|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b153  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [153],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [154]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [152],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [153]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b154|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b155  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [155],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [156]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [154],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [155]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b156|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b157  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [157],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [158]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [156],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [157]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b158|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b159  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [159],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [160]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_13 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [158],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [159]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b160|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b161  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [161],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [162]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [160],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [161]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b162|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b163  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [163],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [164]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [162],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [163]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b164|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b165  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [165],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [166]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [164],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [165]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b166|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b167  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [167],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [168]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [166],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [167]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b168|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b169  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [169],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [170]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [168],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [169]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b16|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b17  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [17],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [18]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_1 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [16],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [17]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b170|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b171  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [171],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [172]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [170],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [171]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b172|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b173  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [173],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [174]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [172],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [173]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b174|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b175  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [175],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [176]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [174],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [175]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b176|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b177  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [177],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [178]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [176],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [177]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b178|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b179  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [179],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [180]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [178],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [179]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b180|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b181  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [181],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [182]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [180],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [181]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b182|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b183  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [183],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [184]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [182],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [183]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b184|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b185  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [185],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [186]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [184],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [185]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b186|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b187  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [187],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [188]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [186],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [187]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b188|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b189  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [189],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [190]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [188],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [189]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b18|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b19  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [19],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [20]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_1 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [18],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [19]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b190|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b191  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [191],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [192]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [190],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [191]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b192|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b193  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [193],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [194]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [192],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [193]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b194|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b195  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [195],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [196]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [194],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [195]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b196|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b197  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [197],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [198]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [196],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [197]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b198|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b199  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [199],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [200]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_13 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [198],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [199]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b1|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b2  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [2],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [3]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [1],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [2]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b200|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b201  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [201],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [202]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [200],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [201]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b202|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b203  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [203],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [204]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [202],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [203]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b204|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b205  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [205],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [206]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [204],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [205]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b206|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b207  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [207],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [208]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [206],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [207]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b208|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b209  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [209],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [210]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [208],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [209]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b20|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b21  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [21],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [22]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_1 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [20],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [21]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b210|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b211  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [211],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [212]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [210],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [211]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b212|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b213  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [213],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [214]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [212],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [213]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b214|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b215  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [215],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [216]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [214],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [215]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b216|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b217  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [217],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [218]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [216],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [217]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b218|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b219  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [219],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [220]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [218],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [219]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b220|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b221  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [221],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [222]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [220],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [221]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b222|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b223  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [223],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [224]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [222],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [223]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b224|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b225  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [225],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [226]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [224],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [225]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b226|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b227  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [227],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [228]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [226],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [227]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b228|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b229  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [229],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [230]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [228],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [229]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b22|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b23  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [23],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [24]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [22],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [23]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b230|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b231  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [231],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [232]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [230],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [231]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b232|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b233  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [233],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [234]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [232],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [233]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b234|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b235  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [235],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [236]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [234],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [235]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b236|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b237  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [237],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [238]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [236],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [237]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b238|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b239  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [239],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [240]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [238],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [239]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b240|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b241  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [241],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [242]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [240],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [241]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b242|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b243  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [243],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [244]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [242],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [243]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b244|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b245  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [245],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [246]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_13 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [244],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [245]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b246|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b247  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [247],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [248]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_13 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [246],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [247]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b248|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b249  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [249],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [250]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_13 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [248],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [249]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b24|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b25  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [25],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [26]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [24],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [25]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b250|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b251  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [251],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [252]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [250],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [251]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b252|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b253  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [253],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [254]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [252],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [253]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b254|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b255  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [255],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [256]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [254],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [255]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b256|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b257  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [257],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [258]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [256],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [257]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b258|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b259  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [259],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [260]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [258],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [259]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b260|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b261  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [261],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [262]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [260],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [261]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b262|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b263  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [263],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [264]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [262],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [263]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b264|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b265  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [265],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [266]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [264],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [265]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b266|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b267  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [267],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [268]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [266],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [267]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b268|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b269  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [269],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [270]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [268],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [269]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b26|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b27  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [27],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [28]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [26],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [27]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b270|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b271  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [271],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [272]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [270],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [271]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b272|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b273  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [273],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [274]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [272],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [273]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b274|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b275  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [275],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [276]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [274],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [275]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b276|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b277  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [277],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [278]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [276],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [277]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b278|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b279  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [279],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [280]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [278],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [279]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b280|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b281  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [281],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [282]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [280],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [281]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b282|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b283  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [283],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [284]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [282],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [283]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b284|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b285  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [285],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [286]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [284],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [285]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b286|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b287  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [287],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [288]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [286],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [287]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b288|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b289  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [289],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [290]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [288],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [289]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b28|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b29  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [29],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [30]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [28],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [29]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b290|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b291  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [291],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [292]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [290],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [291]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b292|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b293  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [293],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [294]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [292],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [293]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b294|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b295  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [295],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [296]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [294],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [295]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b296|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b297  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [297],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [298]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [296],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [297]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b298|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b299  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [299],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [300]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [298],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [299]}));  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b3  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({open_n28428,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [4]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 ),
    .q({open_n28434,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [3]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b300|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b301  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [301],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [302]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [300],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [301]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b302|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b303  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [303],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [304]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [302],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [303]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b304|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b305  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [305],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [306]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [304],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [305]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b306|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b307  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [307],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [308]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [306],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [307]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b308|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b309  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [309],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [310]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [308],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [309]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b30|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b31  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [31],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [32]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [30],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [31]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b310|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b311  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [311],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [312]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [310],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [311]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_LSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b312|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b0  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({jtdi,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [1]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [312],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [0]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b32|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b33  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [33],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [34]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [32],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [33]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b34|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b35  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [35],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [36]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [34],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [35]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b36|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b37  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [37],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [38]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [36],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [37]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b38|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b39  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [39],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [40]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [38],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [39]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b40|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b41  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [41],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [42]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [40],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [41]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b42|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b43  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [43],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [44]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [42],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [43]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b44|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b45  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [45],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [46]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [44],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [45]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b46|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b47  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [47],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [48]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [46],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [47]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b48|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b49  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [49],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [50]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [48],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [49]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b4|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b5  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [5],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [6]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [4],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [5]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b50|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b51  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [51],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [52]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [50],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [51]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b52|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b53  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [53],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [54]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [52],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [53]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b54|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b55  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [55],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [56]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [54],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [55]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b56|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b57  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [57],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [58]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [56],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [57]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b58|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b59  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [59],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [60]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [58],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [59]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b60|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b61  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [61],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [62]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [60],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [61]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b62|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b63  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [63],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [64]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [62],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [63]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b64|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b65  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [65],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [66]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [64],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [65]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b66|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b67  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [67],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [68]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [66],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [67]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b68|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b69  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [69],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [70]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [68],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [69]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b6|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b7  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [7],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [8]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_1 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [6],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [7]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b70|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b71  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [71],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [72]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [70],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [71]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b72|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b73  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [73],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [74]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [72],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [73]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b74|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b75  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [75],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [76]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [74],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [75]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b76|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b77  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [77],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [78]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [76],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [77]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b78|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b79  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [79],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [80]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [78],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [79]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b80|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b81  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [81],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [82]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [80],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [81]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b82|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b83  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [83],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [84]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [82],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [83]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b84|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b85  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [85],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [86]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [84],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [85]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b86|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b87  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [87],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [88]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [86],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [87]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b88|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b89  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [89],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [90]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [88],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [89]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b8|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b9  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [9],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [10]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_1 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [8],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [9]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b90|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b91  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [91],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [92]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [90],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [91]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b92|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b93  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [93],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [94]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [92],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [93]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b94|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b95  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [95],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [96]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [94],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [95]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b96|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b97  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [97],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [98]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [96],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [97]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\register.v(23)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/reg_inst/reg2_b98|cfg_int/wrapper_cfg_inst/reg_inst/reg2_b99  (
    .ce(\cfg_int/wrapper_cfg_inst/shift_0 ),
    .clk(jtck),
    .mi({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [99],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [100]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 ),
    .q({\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [98],\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [99]}));  // D:/td/td/cw\register.v(23)
  // D:/td/td/cw\tap.v(32)
  // D:/td/td/cw\tap.v(32)
  EG_PHY_MSLICE #(
    //.LUT0("(D*A)"),
    //.LUT1("(D*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101000000000),
    .INIT_LUT1(16'b0101010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/jscan_1_r2_reg|cfg_int/wrapper_cfg_inst/tap_inst/jscan_1_r_reg  (
    .a({\cfg_int/wrapper_cfg_inst/tap_inst/jscan_1_r2 ,jscan_1}),
    .clk(jtck),
    .d({\cfg_int/wrapper_cfg_inst/tap_inst/jscan_1_r ,jshift}),
    .mi({\cfg_int/wrapper_cfg_inst/tap_inst/jscan_1_r ,jscan_1}),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 ),
    .f({_al_u3034_o,_al_u3035_o}),
    .q({\cfg_int/wrapper_cfg_inst/tap_inst/jscan_1_r2 ,\cfg_int/wrapper_cfg_inst/tap_inst/jscan_1_r }));  // D:/td/td/cw\tap.v(32)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg  (
    .clk(jtck),
    .mi({open_n29511,1'b0}),
    .sr(jrstn),
    .q({open_n29517,\cfg_int/wrapper_cfg_inst/rst }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_1  (
    .clk(jtck),
    .mi({open_n29537,1'b0}),
    .sr(jrstn),
    .q({open_n29543,\cfg_int/wrapper_cfg_inst/rst_placeOpt_1 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_10  (
    .clk(jtck),
    .mi({open_n29563,1'b0}),
    .sr(jrstn),
    .q({open_n29569,\cfg_int/wrapper_cfg_inst/rst_placeOpt_10 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_11  (
    .clk(jtck),
    .mi({open_n29589,1'b0}),
    .sr(jrstn),
    .q({open_n29595,\cfg_int/wrapper_cfg_inst/rst_placeOpt_11 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_12  (
    .clk(jtck),
    .mi({open_n29615,1'b0}),
    .sr(jrstn),
    .q({open_n29621,\cfg_int/wrapper_cfg_inst/rst_placeOpt_12 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_13  (
    .clk(jtck),
    .mi({open_n29641,1'b0}),
    .sr(jrstn),
    .q({open_n29647,\cfg_int/wrapper_cfg_inst/rst_placeOpt_13 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_14  (
    .clk(jtck),
    .mi({open_n29667,1'b0}),
    .sr(jrstn),
    .q({open_n29673,\cfg_int/wrapper_cfg_inst/rst_placeOpt_14 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_15  (
    .clk(jtck),
    .mi({open_n29693,1'b0}),
    .sr(jrstn),
    .q({open_n29699,\cfg_int/wrapper_cfg_inst/rst_placeOpt_15 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_16  (
    .clk(jtck),
    .mi({open_n29719,1'b0}),
    .sr(jrstn),
    .q({open_n29725,\cfg_int/wrapper_cfg_inst/rst_placeOpt_16 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_17  (
    .clk(jtck),
    .mi({open_n29745,1'b0}),
    .sr(jrstn),
    .q({open_n29751,\cfg_int/wrapper_cfg_inst/rst_placeOpt_17 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_2  (
    .clk(jtck),
    .mi({open_n29771,1'b0}),
    .sr(jrstn),
    .q({open_n29777,\cfg_int/wrapper_cfg_inst/rst_placeOpt_2 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_3  (
    .clk(jtck),
    .mi({open_n29797,1'b0}),
    .sr(jrstn),
    .q({open_n29803,\cfg_int/wrapper_cfg_inst/rst_placeOpt_3 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_4  (
    .clk(jtck),
    .mi({open_n29823,1'b0}),
    .sr(jrstn),
    .q({open_n29829,\cfg_int/wrapper_cfg_inst/rst_placeOpt_4 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_5  (
    .clk(jtck),
    .mi({open_n29849,1'b0}),
    .sr(jrstn),
    .q({open_n29855,\cfg_int/wrapper_cfg_inst/rst_placeOpt_5 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_6  (
    .clk(jtck),
    .mi({open_n29875,1'b0}),
    .sr(jrstn),
    .q({open_n29881,\cfg_int/wrapper_cfg_inst/rst_placeOpt_6 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_7  (
    .clk(jtck),
    .mi({open_n29901,1'b0}),
    .sr(jrstn),
    .q({open_n29907,\cfg_int/wrapper_cfg_inst/rst_placeOpt_7 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_8  (
    .clk(jtck),
    .mi({open_n29927,1'b0}),
    .sr(jrstn),
    .q({open_n29933,\cfg_int/wrapper_cfg_inst/rst_placeOpt_8 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \cfg_int/wrapper_cfg_inst/tap_inst/rst_reg_placeOpt_9  (
    .clk(jtck),
    .mi({open_n29953,1'b0}),
    .sr(jrstn),
    .q({open_n29959,\cfg_int/wrapper_cfg_inst/rst_placeOpt_9 }));  // D:/td/td/cw\tap.v(42)
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P138"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("RESET"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTRSTMUX("INV"),
    .OUTSCLKMUX("CLK"),
    .SRMODE("ASYNC"),
    .TSMUX("0"))
    led_n_reg_DO (
    .ce(n7),
    .do({open_n29998,open_n29999,open_n30000,o_data[0]}),
    .osclk(clock_pad),
    .rst(rst_pad),
    .opad(led));  // __top.v(63)
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \lt0_0|lt0_cin  (
    .a({addr[0],1'b0}),
    .b({1'b0,open_n30012}),
    .clk(clock_pad),
    .mi({addr[0],addr[0]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .fco(lt0_c1),
    .q({\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r }));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_10|lt0_9  (
    .a(addr[10:9]),
    .b(2'b00),
    .fci(lt0_c9),
    .fco(lt0_c11));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_12|lt0_11  (
    .a(addr[12:11]),
    .b(2'b00),
    .fci(lt0_c11),
    .fco(lt0_c13));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_14|lt0_13  (
    .a(addr[14:13]),
    .b(2'b00),
    .fci(lt0_c13),
    .fco(lt0_c15));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_16|lt0_15  (
    .a(addr[16:15]),
    .b(2'b00),
    .fci(lt0_c15),
    .fco(lt0_c17));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_18|lt0_17  (
    .a(addr[18:17]),
    .b(2'b00),
    .fci(lt0_c17),
    .fco(lt0_c19));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_20|lt0_19  (
    .a(addr[20:19]),
    .b(2'b00),
    .fci(lt0_c19),
    .fco(lt0_c21));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_22|lt0_21  (
    .a(addr[22:21]),
    .b(2'b00),
    .fci(lt0_c21),
    .fco(lt0_c23));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_24|lt0_23  (
    .a(addr[24:23]),
    .b(2'b00),
    .fci(lt0_c23),
    .fco(lt0_c25));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_26|lt0_25  (
    .a(addr[26:25]),
    .b(2'b00),
    .fci(lt0_c25),
    .fco(lt0_c27));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_28|lt0_27  (
    .a(addr[28:27]),
    .b(2'b00),
    .fci(lt0_c27),
    .fco(lt0_c29));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_2|lt0_1  (
    .a(addr[2:1]),
    .b(2'b00),
    .fci(lt0_c1),
    .fco(lt0_c3));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_30|lt0_29  (
    .a(addr[30:29]),
    .b(2'b00),
    .fci(lt0_c29),
    .fco(lt0_c31));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_4|lt0_3  (
    .a(addr[4:3]),
    .b(2'b00),
    .fci(lt0_c3),
    .fco(lt0_c5));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_6|lt0_5  (
    .a(addr[6:5]),
    .b(2'b11),
    .fci(lt0_c5),
    .fco(lt0_c7));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_8|lt0_7  (
    .a(addr[8:7]),
    .b(2'b00),
    .fci(lt0_c7),
    .fco(lt0_c9));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_cout|lt0_31  (
    .a({1'b0,addr[31]}),
    .b(2'b10),
    .fci(lt0_c31),
    .f({n0,open_n30410}));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c0_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c0_l  (
    .a({o_data[0],n2[0]}),
    .b({o_data[1],n2[1]}),
    .c({o_data[2],n2[2]}),
    .clk(clock_pad),
    .d({o_data[3],n2[3]}),
    .e({open_n30417,memwrite_cs}),
    .dpram_di(\m/dram_c0_di ),
    .dpram_mode(\m/dram_c0_mode ),
    .dpram_waddr(\m/dram_c0_waddr ),
    .dpram_wclk(\m/dram_c0_wclk ),
    .dpram_we(\m/dram_c0_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c0_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000110),
    .INIT_LUT1(16'b0000000000000110),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c0_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_2 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c0_di [1:0]),
    .dpram_mode(\m/dram_c0_mode ),
    .dpram_waddr(\m/dram_c0_waddr ),
    .dpram_wclk(\m/dram_c0_wclk ),
    .dpram_we(\m/dram_c0_we ),
    .sr(rst_pad),
    .f(i_data[1:0]),
    .q(\t/busarbitration/instruction [1:0]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c0_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c0_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_2 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c0_di [3:2]),
    .dpram_mode(\m/dram_c0_mode ),
    .dpram_waddr(\m/dram_c0_waddr ),
    .dpram_wclk(\m/dram_c0_wclk ),
    .dpram_we(\m/dram_c0_we ),
    .sr(rst_pad),
    .f(i_data[3:2]),
    .q(\t/busarbitration/instruction [3:2]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c1_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c1_l  (
    .a({o_data[4],n2[0]}),
    .b({o_data[5],n2[1]}),
    .c({o_data[6],n2[2]}),
    .clk(clock_pad),
    .d({o_data[7],n2[3]}),
    .e({open_n30442,memwrite_cs}),
    .dpram_di(\m/dram_c1_di ),
    .dpram_mode(\m/dram_c1_mode ),
    .dpram_waddr(\m/dram_c1_waddr ),
    .dpram_wclk(\m/dram_c1_wclk ),
    .dpram_we(\m/dram_c1_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c1_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000110),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c1_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_2 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c1_di [1:0]),
    .dpram_mode(\m/dram_c1_mode ),
    .dpram_waddr(\m/dram_c1_waddr ),
    .dpram_wclk(\m/dram_c1_wclk ),
    .dpram_we(\m/dram_c1_we ),
    .sr(rst_pad),
    .f(i_data[5:4]),
    .q(\t/busarbitration/instruction [5:4]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c1_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c1_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_2 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c1_di [3:2]),
    .dpram_mode(\m/dram_c1_mode ),
    .dpram_waddr(\m/dram_c1_waddr ),
    .dpram_wclk(\m/dram_c1_wclk ),
    .dpram_we(\m/dram_c1_we ),
    .sr(rst_pad),
    .f(i_data[7:6]),
    .q(\t/busarbitration/instruction [7:6]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c2_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c2_l  (
    .a({o_data[8],n2[0]}),
    .b({o_data[9],n2[1]}),
    .c({o_data[10],n2[2]}),
    .clk(clock_pad),
    .d({o_data[11],n2[3]}),
    .e({open_n30467,memwrite_cs}),
    .dpram_di(\m/dram_c2_di ),
    .dpram_mode(\m/dram_c2_mode ),
    .dpram_waddr(\m/dram_c2_waddr ),
    .dpram_wclk(\m/dram_c2_wclk ),
    .dpram_we(\m/dram_c2_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c2_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c2_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_2 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c2_di [1:0]),
    .dpram_mode(\m/dram_c2_mode ),
    .dpram_waddr(\m/dram_c2_waddr ),
    .dpram_wclk(\m/dram_c2_wclk ),
    .dpram_we(\m/dram_c2_we ),
    .sr(rst_pad),
    .f(i_data[9:8]),
    .q(\t/busarbitration/instruction [9:8]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c2_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c2_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_2 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c2_di [3:2]),
    .dpram_mode(\m/dram_c2_mode ),
    .dpram_waddr(\m/dram_c2_waddr ),
    .dpram_wclk(\m/dram_c2_wclk ),
    .dpram_we(\m/dram_c2_we ),
    .sr(rst_pad),
    .f(i_data[11:10]),
    .q(\t/busarbitration/instruction [11:10]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c3_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c3_l  (
    .a({o_data[12],n2[0]}),
    .b({o_data[13],n2[1]}),
    .c({o_data[14],n2[2]}),
    .clk(clock_pad),
    .d({o_data[15],n2[3]}),
    .e({open_n30492,memwrite_cs}),
    .dpram_di(\m/dram_c3_di ),
    .dpram_mode(\m/dram_c3_mode ),
    .dpram_waddr(\m/dram_c3_waddr ),
    .dpram_wclk(\m/dram_c3_wclk ),
    .dpram_we(\m/dram_c3_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c3_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000110),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c3_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_5 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c3_di [1:0]),
    .dpram_mode(\m/dram_c3_mode ),
    .dpram_waddr(\m/dram_c3_waddr ),
    .dpram_wclk(\m/dram_c3_wclk ),
    .dpram_we(\m/dram_c3_we ),
    .sr(rst_pad),
    .f(i_data[13:12]),
    .q(\t/busarbitration/instruction [13:12]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c3_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000110),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c3_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_5 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c3_di [3:2]),
    .dpram_mode(\m/dram_c3_mode ),
    .dpram_waddr(\m/dram_c3_waddr ),
    .dpram_wclk(\m/dram_c3_wclk ),
    .dpram_we(\m/dram_c3_we ),
    .sr(rst_pad),
    .f(i_data[15:14]),
    .q(\t/busarbitration/instruction [15:14]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c4_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c4_l  (
    .a({o_data[16],n2[0]}),
    .b({o_data[17],n2[1]}),
    .c({o_data[18],n2[2]}),
    .clk(clock_pad),
    .d({o_data[19],n2[3]}),
    .e({open_n30517,memwrite_cs}),
    .dpram_di(\m/dram_c4_di ),
    .dpram_mode(\m/dram_c4_mode ),
    .dpram_waddr(\m/dram_c4_waddr ),
    .dpram_wclk(\m/dram_c4_wclk ),
    .dpram_we(\m/dram_c4_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c4_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c4_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_5 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c4_di [1:0]),
    .dpram_mode(\m/dram_c4_mode ),
    .dpram_waddr(\m/dram_c4_waddr ),
    .dpram_wclk(\m/dram_c4_wclk ),
    .dpram_we(\m/dram_c4_we ),
    .sr(rst_pad),
    .f(i_data[17:16]),
    .q(\t/busarbitration/instruction [17:16]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c4_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c4_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_5 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c4_di [3:2]),
    .dpram_mode(\m/dram_c4_mode ),
    .dpram_waddr(\m/dram_c4_waddr ),
    .dpram_wclk(\m/dram_c4_wclk ),
    .dpram_we(\m/dram_c4_we ),
    .sr(rst_pad),
    .f(i_data[19:18]),
    .q(\t/busarbitration/instruction [19:18]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c5_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c5_l  (
    .a({o_data[20],n2[0]}),
    .b({o_data[21],n2[1]}),
    .c({o_data[22],n2[2]}),
    .clk(clock_pad),
    .d({o_data[23],n2[3]}),
    .e({open_n30542,memwrite_cs}),
    .dpram_di(\m/dram_c5_di ),
    .dpram_mode(\m/dram_c5_mode ),
    .dpram_waddr(\m/dram_c5_waddr ),
    .dpram_wclk(\m/dram_c5_wclk ),
    .dpram_we(\m/dram_c5_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c5_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c5_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_5 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c5_di [1:0]),
    .dpram_mode(\m/dram_c5_mode ),
    .dpram_waddr(\m/dram_c5_waddr ),
    .dpram_wclk(\m/dram_c5_wclk ),
    .dpram_we(\m/dram_c5_we ),
    .sr(rst_pad),
    .f(i_data[21:20]),
    .q(\t/busarbitration/instruction [21:20]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c5_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c5_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_5 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c5_di [3:2]),
    .dpram_mode(\m/dram_c5_mode ),
    .dpram_waddr(\m/dram_c5_waddr ),
    .dpram_wclk(\m/dram_c5_wclk ),
    .dpram_we(\m/dram_c5_we ),
    .sr(rst_pad),
    .f(i_data[23:22]),
    .q(\t/busarbitration/instruction [23:22]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c6_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c6_l  (
    .a({o_data[24],n2[0]}),
    .b({o_data[25],n2[1]}),
    .c({o_data[26],n2[2]}),
    .clk(clock_pad),
    .d({o_data[27],n2[3]}),
    .e({open_n30567,memwrite_cs}),
    .dpram_di(\m/dram_c6_di ),
    .dpram_mode(\m/dram_c6_mode ),
    .dpram_waddr(\m/dram_c6_waddr ),
    .dpram_wclk(\m/dram_c6_wclk ),
    .dpram_we(\m/dram_c6_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c6_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c6_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_5 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c6_di [1:0]),
    .dpram_mode(\m/dram_c6_mode ),
    .dpram_waddr(\m/dram_c6_waddr ),
    .dpram_wclk(\m/dram_c6_wclk ),
    .dpram_we(\m/dram_c6_we ),
    .sr(rst_pad),
    .f(i_data[25:24]),
    .q(\t/busarbitration/instruction [25:24]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c6_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c6_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_5 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c6_di [3:2]),
    .dpram_mode(\m/dram_c6_mode ),
    .dpram_waddr(\m/dram_c6_waddr ),
    .dpram_wclk(\m/dram_c6_wclk ),
    .dpram_we(\m/dram_c6_we ),
    .sr(rst_pad),
    .f(i_data[27:26]),
    .q(\t/busarbitration/instruction [27:26]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c7_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c7_l  (
    .a({o_data[28],n2[0]}),
    .b({o_data[29],n2[1]}),
    .c({o_data[30],n2[2]}),
    .clk(clock_pad),
    .d({o_data[31],n2[3]}),
    .e({open_n30592,memwrite_cs}),
    .dpram_di(\m/dram_c7_di ),
    .dpram_mode(\m/dram_c7_mode ),
    .dpram_waddr(\m/dram_c7_waddr ),
    .dpram_wclk(\m/dram_c7_wclk ),
    .dpram_we(\m/dram_c7_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c7_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c7_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_5 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c7_di [1:0]),
    .dpram_mode(\m/dram_c7_mode ),
    .dpram_waddr(\m/dram_c7_waddr ),
    .dpram_wclk(\m/dram_c7_wclk ),
    .dpram_we(\m/dram_c7_we ),
    .sr(rst_pad),
    .f(i_data[29:28]),
    .q(\t/busarbitration/instruction [29:28]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c7_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000110),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c7_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3_placeOpt_5 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c7_di [3:2]),
    .dpram_mode(\m/dram_c7_mode ),
    .dpram_waddr(\m/dram_c7_waddr ),
    .dpram_wclk(\m/dram_c7_wclk ),
    .dpram_we(\m/dram_c7_we ),
    .sr(rst_pad),
    .f(i_data[31:30]),
    .q(\t/busarbitration/instruction [31:30]));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u11_al_u2928  (
    .a({\t/a/EX_A [13],\t/a/EX_A [11]}),
    .b({\t/a/EX_A [14],\t/a/EX_A [12]}),
    .c(2'b00),
    .d({\t/a/EX_B [13],\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/EX_B [14],\t/a/EX_B [12]}),
    .fci(\t/a/alu/add0/c11 ),
    .f({\t/a/alu/n5 [13],\t/a/alu/n5 [11]}),
    .fco(\t/a/alu/add0/c15 ),
    .fx({\t/a/alu/n5 [14],\t/a/alu/n5 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u15_al_u2929  (
    .a({\t/a/EX_A [17],\t/a/EX_A [15]}),
    .b({\t/a/EX_A [18],\t/a/EX_A [16]}),
    .c(2'b00),
    .d({\t/a/EX_B [17],\t/a/EX_B [15]}),
    .e({\t/a/EX_B [18],\t/a/EX_B [16]}),
    .fci(\t/a/alu/add0/c15 ),
    .f({\t/a/alu/n5 [17],\t/a/alu/n5 [15]}),
    .fco(\t/a/alu/add0/c19 ),
    .fx({\t/a/alu/n5 [18],\t/a/alu/n5 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u19_al_u2930  (
    .a({\t/a/EX_A [21],\t/a/EX_A [19]}),
    .b({\t/a/EX_A [22],\t/a/EX_A [20]}),
    .c(2'b00),
    .d({\t/a/EX_B [21],\t/a/EX_B [19]}),
    .e({\t/a/EX_B [22],\t/a/EX_B [20]}),
    .fci(\t/a/alu/add0/c19 ),
    .f({\t/a/alu/n5 [21],\t/a/alu/n5 [19]}),
    .fco(\t/a/alu/add0/c23 ),
    .fx({\t/a/alu/n5 [22],\t/a/alu/n5 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u23_al_u2931  (
    .a({\t/a/EX_A [25],\t/a/EX_A [23]}),
    .b({\t/a/EX_A [26],\t/a/EX_A [24]}),
    .c(2'b00),
    .d({\t/a/EX_B [25],\t/a/EX_B [23]}),
    .e({\t/a/EX_B [26],\t/a/EX_B [24]}),
    .fci(\t/a/alu/add0/c23 ),
    .f({\t/a/alu/n5 [25],\t/a/alu/n5 [23]}),
    .fco(\t/a/alu/add0/c27 ),
    .fx({\t/a/alu/n5 [26],\t/a/alu/n5 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u27_al_u2932  (
    .a({\t/a/EX_A [29],\t/a/EX_A [27]}),
    .b({\t/a/EX_A [30],\t/a/EX_A [28]}),
    .c(2'b00),
    .d({\t/a/EX_B [29],\t/a/EX_B [27]}),
    .e({\t/a/EX_B [30],\t/a/EX_B [28]}),
    .fci(\t/a/alu/add0/c27 ),
    .f({\t/a/alu/n5 [29],\t/a/alu/n5 [27]}),
    .fco(\t/a/alu/add0/c31 ),
    .fx({\t/a/alu/n5 [30],\t/a/alu/n5 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u31_al_u2933  (
    .a({open_n30706,\t/a/EX_A [31]}),
    .c(2'b00),
    .d({open_n30711,\t/a/EX_B [31]}),
    .fci(\t/a/alu/add0/c31 ),
    .f({open_n30728,\t/a/alu/n5 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u3_al_u2926  (
    .a({\t/a/EX_A [5],\t/a/EX_A [3]}),
    .b({\t/a/EX_A [6],\t/a/EX_A [4]}),
    .c(2'b00),
    .d({\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_1 }),
    .e({\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/add0/c3 ),
    .f({\t/a/alu/n5 [5],\t/a/alu/n5 [3]}),
    .fco(\t/a/alu/add0/c7 ),
    .fx({\t/a/alu/n5 [6],\t/a/alu/n5 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u7_al_u2927  (
    .a({\t/a/EX_A [9],\t/a/EX_A [7]}),
    .b({\t/a/EX_A [10],\t/a/EX_A [8]}),
    .c(2'b00),
    .d({\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/add0/c7 ),
    .f({\t/a/alu/n5 [9],\t/a/alu/n5 [7]}),
    .fco(\t/a/alu/add0/c11 ),
    .fx({\t/a/alu/n5 [10],\t/a/alu/n5 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/ucin_al_u2925  (
    .a({\t/a/EX_A [1],1'b0}),
    .b({\t/a/EX_A [2],\t/a/EX_A [0]}),
    .c(2'b00),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,1'b1}),
    .e({\t/a/EX_B [2],\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({\t/a/alu/n5 [1],open_n30787}),
    .fco(\t/a/alu/add0/c3 ),
    .fx({\t/a/alu/n5 [2],\t/a/alu/n5 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_0|t/a/alu/lt0_cin  (
    .a({\t/a/EX_A [0],1'b0}),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,open_n30790}),
    .fco(\t/a/alu/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_10|t/a/alu/lt0_9  (
    .a(\t/a/EX_A [10:9]),
    .b({\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/lt0_c9 ),
    .fco(\t/a/alu/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_12|t/a/alu/lt0_11  (
    .a(\t/a/EX_A [12:11]),
    .b({\t/a/EX_B [12],\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/lt0_c11 ),
    .fco(\t/a/alu/lt0_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_14|t/a/alu/lt0_13  (
    .a(\t/a/EX_A [14:13]),
    .b(\t/a/EX_B [14:13]),
    .fci(\t/a/alu/lt0_c13 ),
    .fco(\t/a/alu/lt0_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_16|t/a/alu/lt0_15  (
    .a(\t/a/EX_A [16:15]),
    .b(\t/a/EX_B [16:15]),
    .fci(\t/a/alu/lt0_c15 ),
    .fco(\t/a/alu/lt0_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_18|t/a/alu/lt0_17  (
    .a(\t/a/EX_A [18:17]),
    .b(\t/a/EX_B [18:17]),
    .fci(\t/a/alu/lt0_c17 ),
    .fco(\t/a/alu/lt0_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_20|t/a/alu/lt0_19  (
    .a(\t/a/EX_A [20:19]),
    .b(\t/a/EX_B [20:19]),
    .fci(\t/a/alu/lt0_c19 ),
    .fco(\t/a/alu/lt0_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_22|t/a/alu/lt0_21  (
    .a(\t/a/EX_A [22:21]),
    .b(\t/a/EX_B [22:21]),
    .fci(\t/a/alu/lt0_c21 ),
    .fco(\t/a/alu/lt0_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_24|t/a/alu/lt0_23  (
    .a(\t/a/EX_A [24:23]),
    .b(\t/a/EX_B [24:23]),
    .fci(\t/a/alu/lt0_c23 ),
    .fco(\t/a/alu/lt0_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_26|t/a/alu/lt0_25  (
    .a(\t/a/EX_A [26:25]),
    .b(\t/a/EX_B [26:25]),
    .fci(\t/a/alu/lt0_c25 ),
    .fco(\t/a/alu/lt0_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_28|t/a/alu/lt0_27  (
    .a(\t/a/EX_A [28:27]),
    .b(\t/a/EX_B [28:27]),
    .fci(\t/a/alu/lt0_c27 ),
    .fco(\t/a/alu/lt0_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_2|t/a/alu/lt0_1  (
    .a(\t/a/EX_A [2:1]),
    .b({\t/a/EX_B [2],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/lt0_c1 ),
    .fco(\t/a/alu/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_30|t/a/alu/lt0_29  (
    .a(\t/a/EX_A [30:29]),
    .b(\t/a/EX_B [30:29]),
    .fci(\t/a/alu/lt0_c29 ),
    .fco(\t/a/alu/lt0_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_4|t/a/alu/lt0_3  (
    .a(\t/a/EX_A [4:3]),
    .b({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_3 }),
    .fci(\t/a/alu/lt0_c3 ),
    .fco(\t/a/alu/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_6|t/a/alu/lt0_5  (
    .a(\t/a/EX_A [6:5]),
    .b({\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/lt0_c5 ),
    .fco(\t/a/alu/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_8|t/a/alu/lt0_7  (
    .a(\t/a/EX_A [8:7]),
    .b({\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/lt0_c7 ),
    .fco(\t/a/alu/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_cout|t/a/alu/lt0_31  (
    .a({1'b0,\t/a/EX_A [31]}),
    .b({1'b1,\t/a/EX_B [31]}),
    .fci(\t/a/alu/lt0_c31 ),
    .f({\t/a/alu/n8 ,open_n31194}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u11_al_u2937  (
    .a({\t/a/EX_A [13],\t/a/EX_A [11]}),
    .b({\t/a/EX_A [14],\t/a/EX_A [12]}),
    .c(2'b11),
    .d({\t/a/EX_B [13],\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/EX_B [14],\t/a/EX_B [12]}),
    .fci(\t/a/alu/sub0/c11 ),
    .f({\t/a/alu/n6 [13],\t/a/alu/n6 [11]}),
    .fco(\t/a/alu/sub0/c15 ),
    .fx({\t/a/alu/n6 [14],\t/a/alu/n6 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u15_al_u2938  (
    .a({\t/a/EX_A [17],\t/a/EX_A [15]}),
    .b({\t/a/EX_A [18],\t/a/EX_A [16]}),
    .c(2'b11),
    .d({\t/a/EX_B [17],\t/a/EX_B [15]}),
    .e({\t/a/EX_B [18],\t/a/EX_B [16]}),
    .fci(\t/a/alu/sub0/c15 ),
    .f({\t/a/alu/n6 [17],\t/a/alu/n6 [15]}),
    .fco(\t/a/alu/sub0/c19 ),
    .fx({\t/a/alu/n6 [18],\t/a/alu/n6 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u19_al_u2939  (
    .a({\t/a/EX_A [21],\t/a/EX_A [19]}),
    .b({\t/a/EX_A [22],\t/a/EX_A [20]}),
    .c(2'b11),
    .d({\t/a/EX_B [21],\t/a/EX_B [19]}),
    .e({\t/a/EX_B [22],\t/a/EX_B [20]}),
    .fci(\t/a/alu/sub0/c19 ),
    .f({\t/a/alu/n6 [21],\t/a/alu/n6 [19]}),
    .fco(\t/a/alu/sub0/c23 ),
    .fx({\t/a/alu/n6 [22],\t/a/alu/n6 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u23_al_u2940  (
    .a({\t/a/EX_A [25],\t/a/EX_A [23]}),
    .b({\t/a/EX_A [26],\t/a/EX_A [24]}),
    .c(2'b11),
    .d({\t/a/EX_B [25],\t/a/EX_B [23]}),
    .e({\t/a/EX_B [26],\t/a/EX_B [24]}),
    .fci(\t/a/alu/sub0/c23 ),
    .f({\t/a/alu/n6 [25],\t/a/alu/n6 [23]}),
    .fco(\t/a/alu/sub0/c27 ),
    .fx({\t/a/alu/n6 [26],\t/a/alu/n6 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u27_al_u2941  (
    .a({\t/a/EX_A [29],\t/a/EX_A [27]}),
    .b({\t/a/EX_A [30],\t/a/EX_A [28]}),
    .c(2'b11),
    .d({\t/a/EX_B [29],\t/a/EX_B [27]}),
    .e({\t/a/EX_B [30],\t/a/EX_B [28]}),
    .fci(\t/a/alu/sub0/c27 ),
    .f({\t/a/alu/n6 [29],\t/a/alu/n6 [27]}),
    .fco(\t/a/alu/sub0/c31 ),
    .fx({\t/a/alu/n6 [30],\t/a/alu/n6 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u31_al_u2942  (
    .a({open_n31290,\t/a/EX_A [31]}),
    .c(2'b11),
    .d({open_n31295,\t/a/EX_B [31]}),
    .fci(\t/a/alu/sub0/c31 ),
    .f({open_n31312,\t/a/alu/n6 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u3_al_u2935  (
    .a({\t/a/EX_A [5],\t/a/EX_A [3]}),
    .b({\t/a/EX_A [6],\t/a/EX_A [4]}),
    .c(2'b11),
    .d({\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o_placeOpt_3 }),
    .e({\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/sub0/c3 ),
    .f({\t/a/alu/n6 [5],\t/a/alu/n6 [3]}),
    .fco(\t/a/alu/sub0/c7 ),
    .fx({\t/a/alu/n6 [6],\t/a/alu/n6 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u7_al_u2936  (
    .a({\t/a/EX_A [9],\t/a/EX_A [7]}),
    .b({\t/a/EX_A [10],\t/a/EX_A [8]}),
    .c(2'b11),
    .d({\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/sub0/c7 ),
    .f({\t/a/alu/n6 [9],\t/a/alu/n6 [7]}),
    .fco(\t/a/alu/sub0/c11 ),
    .fx({\t/a/alu/n6 [10],\t/a/alu/n6 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/ucin_al_u2934  (
    .a({\t/a/EX_A [1],1'b0}),
    .b({\t/a/EX_A [2],\t/a/EX_A [0]}),
    .c(2'b11),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,1'b1}),
    .e({\t/a/EX_B [2],\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({\t/a/alu/n6 [1],open_n31371}),
    .fco(\t/a/alu/sub0/c3 ),
    .fx({\t/a/alu/n6 [2],\t/a/alu/n6 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u11_al_u2946  (
    .a({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .b({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [13],\t/a/ID_jump_regdat1 [11]}),
    .e({\t/a/ID_jump_regdat1 [14],\t/a/ID_jump_regdat1 [12]}),
    .fci(\t/a/condition/add0/c11 ),
    .f({\t/a/condition/n5 [13],\t/a/condition/n5 [11]}),
    .fco(\t/a/condition/add0/c15 ),
    .fx({\t/a/condition/n5 [14],\t/a/condition/n5 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u15_al_u2947  (
    .a({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .b({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [17],\t/a/ID_jump_regdat1 [15]}),
    .e({\t/a/ID_jump_regdat1 [18],\t/a/ID_jump_regdat1 [16]}),
    .fci(\t/a/condition/add0/c15 ),
    .f({\t/a/condition/n5 [17],\t/a/condition/n5 [15]}),
    .fco(\t/a/condition/add0/c19 ),
    .fx({\t/a/condition/n5 [18],\t/a/condition/n5 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u19_al_u2948  (
    .a({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .b({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [21],\t/a/ID_jump_regdat1 [19]}),
    .e({\t/a/ID_jump_regdat1 [22],\t/a/ID_jump_regdat1 [20]}),
    .fci(\t/a/condition/add0/c19 ),
    .f({\t/a/condition/n5 [21],\t/a/condition/n5 [19]}),
    .fco(\t/a/condition/add0/c23 ),
    .fx({\t/a/condition/n5 [22],\t/a/condition/n5 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u23_al_u2949  (
    .a({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .b({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [25],\t/a/ID_jump_regdat1 [23]}),
    .e({\t/a/ID_jump_regdat1 [26],\t/a/ID_jump_regdat1 [24]}),
    .fci(\t/a/condition/add0/c23 ),
    .f({\t/a/condition/n5 [25],\t/a/condition/n5 [23]}),
    .fco(\t/a/condition/add0/c27 ),
    .fx({\t/a/condition/n5 [26],\t/a/condition/n5 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u27_al_u2950  (
    .a({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .b({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [29],\t/a/ID_jump_regdat1 [27]}),
    .e({\t/a/ID_jump_regdat1 [30],\t/a/ID_jump_regdat1 [28]}),
    .fci(\t/a/condition/add0/c27 ),
    .f({\t/a/condition/n5 [29],\t/a/condition/n5 [27]}),
    .fco(\t/a/condition/add0/c31 ),
    .fx({\t/a/condition/n5 [30],\t/a/condition/n5 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u31_al_u2951  (
    .a({open_n31464,\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({open_n31469,\t/a/ID_jump_regdat1 [31]}),
    .fci(\t/a/condition/add0/c31 ),
    .f({open_n31486,\t/a/condition/n5 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u3_al_u2944  (
    .a({\t/a/ID_fun7 [0],\t/a/ID_rs2 [3]}),
    .b({\t/a/ID_fun7 [1],\t/a/ID_rs2 [4]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [5],\t/a/ID_jump_regdat1 [3]}),
    .e({\t/a/ID_jump_regdat1 [6],\t/a/ID_jump_regdat1 [4]}),
    .fci(\t/a/condition/add0/c3 ),
    .f({\t/a/condition/n5 [5],\t/a/condition/n5 [3]}),
    .fco(\t/a/condition/add0/c7 ),
    .fx({\t/a/condition/n5 [6],\t/a/condition/n5 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u7_al_u2945  (
    .a({\t/a/ID_fun7 [4],\t/a/ID_fun7 [2]}),
    .b({\t/a/ID_fun7 [5],\t/a/ID_fun7 [3]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [9],\t/a/ID_jump_regdat1 [7]}),
    .e({\t/a/ID_jump_regdat1 [10],\t/a/ID_jump_regdat1 [8]}),
    .fci(\t/a/condition/add0/c7 ),
    .f({\t/a/condition/n5 [9],\t/a/condition/n5 [7]}),
    .fco(\t/a/condition/add0/c11 ),
    .fx({\t/a/condition/n5 [10],\t/a/condition/n5 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/ucin_al_u2943  (
    .a({\t/a/ID_rs2$1$_placeOpt_9 ,1'b0}),
    .b({\t/a/ID_rs2$2$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_15 }),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [1],1'b1}),
    .e({\t/a/ID_jump_regdat1 [2],\t/a/ID_jump_regdat1 [0]}),
    .f({\t/a/condition/n5 [1],open_n31545}),
    .fco(\t/a/condition/add0/c3 ),
    .fx({\t/a/condition/n5 [2],open_n31546}));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_0|t/a/condition/lt0_cin  (
    .a({\t/a/ID_jump_regdat1 [0],1'b0}),
    .b({\t/a/ID_jump_regdat2 [0],open_n31549}),
    .fco(\t/a/condition/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_10|t/a/condition/lt0_9  (
    .a(\t/a/ID_jump_regdat1 [10:9]),
    .b(\t/a/ID_jump_regdat2 [10:9]),
    .fci(\t/a/condition/lt0_c9 ),
    .fco(\t/a/condition/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_12|t/a/condition/lt0_11  (
    .a(\t/a/ID_jump_regdat1 [12:11]),
    .b(\t/a/ID_jump_regdat2 [12:11]),
    .fci(\t/a/condition/lt0_c11 ),
    .fco(\t/a/condition/lt0_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_14|t/a/condition/lt0_13  (
    .a(\t/a/ID_jump_regdat1 [14:13]),
    .b(\t/a/ID_jump_regdat2 [14:13]),
    .fci(\t/a/condition/lt0_c13 ),
    .fco(\t/a/condition/lt0_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_16|t/a/condition/lt0_15  (
    .a(\t/a/ID_jump_regdat1 [16:15]),
    .b(\t/a/ID_jump_regdat2 [16:15]),
    .fci(\t/a/condition/lt0_c15 ),
    .fco(\t/a/condition/lt0_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_18|t/a/condition/lt0_17  (
    .a(\t/a/ID_jump_regdat1 [18:17]),
    .b(\t/a/ID_jump_regdat2 [18:17]),
    .fci(\t/a/condition/lt0_c17 ),
    .fco(\t/a/condition/lt0_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_20|t/a/condition/lt0_19  (
    .a(\t/a/ID_jump_regdat1 [20:19]),
    .b(\t/a/ID_jump_regdat2 [20:19]),
    .fci(\t/a/condition/lt0_c19 ),
    .fco(\t/a/condition/lt0_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_22|t/a/condition/lt0_21  (
    .a(\t/a/ID_jump_regdat1 [22:21]),
    .b(\t/a/ID_jump_regdat2 [22:21]),
    .fci(\t/a/condition/lt0_c21 ),
    .fco(\t/a/condition/lt0_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_24|t/a/condition/lt0_23  (
    .a(\t/a/ID_jump_regdat1 [24:23]),
    .b(\t/a/ID_jump_regdat2 [24:23]),
    .fci(\t/a/condition/lt0_c23 ),
    .fco(\t/a/condition/lt0_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_26|t/a/condition/lt0_25  (
    .a(\t/a/ID_jump_regdat1 [26:25]),
    .b(\t/a/ID_jump_regdat2 [26:25]),
    .fci(\t/a/condition/lt0_c25 ),
    .fco(\t/a/condition/lt0_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_28|t/a/condition/lt0_27  (
    .a(\t/a/ID_jump_regdat1 [28:27]),
    .b(\t/a/ID_jump_regdat2 [28:27]),
    .fci(\t/a/condition/lt0_c27 ),
    .fco(\t/a/condition/lt0_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_2|t/a/condition/lt0_1  (
    .a(\t/a/ID_jump_regdat1 [2:1]),
    .b(\t/a/ID_jump_regdat2 [2:1]),
    .fci(\t/a/condition/lt0_c1 ),
    .fco(\t/a/condition/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_30|t/a/condition/lt0_29  (
    .a(\t/a/ID_jump_regdat1 [30:29]),
    .b(\t/a/ID_jump_regdat2 [30:29]),
    .fci(\t/a/condition/lt0_c29 ),
    .fco(\t/a/condition/lt0_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_4|t/a/condition/lt0_3  (
    .a(\t/a/ID_jump_regdat1 [4:3]),
    .b(\t/a/ID_jump_regdat2 [4:3]),
    .fci(\t/a/condition/lt0_c3 ),
    .fco(\t/a/condition/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_6|t/a/condition/lt0_5  (
    .a(\t/a/ID_jump_regdat1 [6:5]),
    .b(\t/a/ID_jump_regdat2 [6:5]),
    .fci(\t/a/condition/lt0_c5 ),
    .fco(\t/a/condition/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_8|t/a/condition/lt0_7  (
    .a(\t/a/ID_jump_regdat1 [8:7]),
    .b(\t/a/ID_jump_regdat2 [8:7]),
    .fci(\t/a/condition/lt0_c7 ),
    .fco(\t/a/condition/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_cout|t/a/condition/lt0_31  (
    .a({1'b0,\t/a/ID_jump_regdat1 [31]}),
    .b({1'b1,\t/a/ID_jump_regdat2 [31]}),
    .fci(\t/a/condition/lt0_c31 ),
    .f({\t/a/condition/n9 ,open_n31953}));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_0|t/a/condition/lt1_cin  (
    .a({\t/a/ID_jump_regdat1 [0],1'b0}),
    .b({\t/a/ID_jump_regdat2 [0],open_n31959}),
    .fco(\t/a/condition/lt1_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_10|t/a/condition/lt1_9  (
    .a(\t/a/ID_jump_regdat1 [10:9]),
    .b(\t/a/ID_jump_regdat2 [10:9]),
    .fci(\t/a/condition/lt1_c9 ),
    .fco(\t/a/condition/lt1_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_12|t/a/condition/lt1_11  (
    .a(\t/a/ID_jump_regdat1 [12:11]),
    .b(\t/a/ID_jump_regdat2 [12:11]),
    .fci(\t/a/condition/lt1_c11 ),
    .fco(\t/a/condition/lt1_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_14|t/a/condition/lt1_13  (
    .a(\t/a/ID_jump_regdat1 [14:13]),
    .b(\t/a/ID_jump_regdat2 [14:13]),
    .fci(\t/a/condition/lt1_c13 ),
    .fco(\t/a/condition/lt1_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_16|t/a/condition/lt1_15  (
    .a(\t/a/ID_jump_regdat1 [16:15]),
    .b(\t/a/ID_jump_regdat2 [16:15]),
    .fci(\t/a/condition/lt1_c15 ),
    .fco(\t/a/condition/lt1_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_18|t/a/condition/lt1_17  (
    .a(\t/a/ID_jump_regdat1 [18:17]),
    .b(\t/a/ID_jump_regdat2 [18:17]),
    .fci(\t/a/condition/lt1_c17 ),
    .fco(\t/a/condition/lt1_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_20|t/a/condition/lt1_19  (
    .a(\t/a/ID_jump_regdat1 [20:19]),
    .b(\t/a/ID_jump_regdat2 [20:19]),
    .fci(\t/a/condition/lt1_c19 ),
    .fco(\t/a/condition/lt1_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_22|t/a/condition/lt1_21  (
    .a(\t/a/ID_jump_regdat1 [22:21]),
    .b(\t/a/ID_jump_regdat2 [22:21]),
    .fci(\t/a/condition/lt1_c21 ),
    .fco(\t/a/condition/lt1_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_24|t/a/condition/lt1_23  (
    .a(\t/a/ID_jump_regdat1 [24:23]),
    .b(\t/a/ID_jump_regdat2 [24:23]),
    .fci(\t/a/condition/lt1_c23 ),
    .fco(\t/a/condition/lt1_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_26|t/a/condition/lt1_25  (
    .a(\t/a/ID_jump_regdat1 [26:25]),
    .b(\t/a/ID_jump_regdat2 [26:25]),
    .fci(\t/a/condition/lt1_c25 ),
    .fco(\t/a/condition/lt1_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_28|t/a/condition/lt1_27  (
    .a(\t/a/ID_jump_regdat1 [28:27]),
    .b(\t/a/ID_jump_regdat2 [28:27]),
    .fci(\t/a/condition/lt1_c27 ),
    .fco(\t/a/condition/lt1_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_2|t/a/condition/lt1_1  (
    .a(\t/a/ID_jump_regdat1 [2:1]),
    .b(\t/a/ID_jump_regdat2 [2:1]),
    .fci(\t/a/condition/lt1_c1 ),
    .fco(\t/a/condition/lt1_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_30|t/a/condition/lt1_29  (
    .a(\t/a/ID_jump_regdat1 [30:29]),
    .b(\t/a/ID_jump_regdat2 [30:29]),
    .fci(\t/a/condition/lt1_c29 ),
    .fco(\t/a/condition/lt1_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_4|t/a/condition/lt1_3  (
    .a(\t/a/ID_jump_regdat1 [4:3]),
    .b(\t/a/ID_jump_regdat2 [4:3]),
    .fci(\t/a/condition/lt1_c3 ),
    .fco(\t/a/condition/lt1_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_6|t/a/condition/lt1_5  (
    .a(\t/a/ID_jump_regdat1 [6:5]),
    .b(\t/a/ID_jump_regdat2 [6:5]),
    .fci(\t/a/condition/lt1_c5 ),
    .fco(\t/a/condition/lt1_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_8|t/a/condition/lt1_7  (
    .a(\t/a/ID_jump_regdat1 [8:7]),
    .b(\t/a/ID_jump_regdat2 [8:7]),
    .fci(\t/a/condition/lt1_c7 ),
    .fco(\t/a/condition/lt1_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_cout_al_u2977  (
    .a({open_n32345,1'b0}),
    .b({open_n32346,1'b1}),
    .fci(\t/a/condition/lt1_c31 ),
    .f({open_n32365,\t/a/condition/n10 }));
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~A*~B*~D+C*~A*~B*~D+~C*~A*B*~D+C*~A*B*~D+~C*~A*~B*D+C*~A*~B*D+~C*A*~B*D+C*A*~B*D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D"),
    //.LUTG0("~C*~A*B*~D+C*~A*B*~D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111101010101),
    .INIT_LUTF1(16'b0111011101110111),
    .INIT_LUTG0(16'b1100110001000100),
    .INIT_LUTG1(16'b0000000001110111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg0_b1|t/a/mem_wb/reg2_b1  (
    .a({_al_u1984_o,\t/a/MEM_rd [4]}),
    .b({\t/a/EX_rs2 [1],\t/a/EX_rs2 [1]}),
    .clk(clock_pad),
    .d({\t/a/EX_rd [1],\t/a/EX_rs2 [4]}),
    .e({\t/a/aluin/n12_lutinv ,\t/a/MEM_rd [1]}),
    .mi({\t/a/EX_rd [1],\t/a/MEM_rd [1]}),
    .sr(rst_pad),
    .f({_al_u2073_o,_al_u1969_o}),
    .q({\t/a/MEM_rd [1],\t/a/WB_rd [1]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*A*~C*D+B*A*~C*D+~B*A*C*D+B*A*C*D"),
    //.LUTF1("~B*~C*~A*~D+B*~C*~A*~D+~B*C*~A*~D+B*C*~A*~D+~B*~C*A*~D+B*~C*A*~D+~B*~C*~A*D+B*~C*~A*D+~B*C*~A*D+B*C*~A*D+~B*~C*A*D+B*~C*A*D"),
    //.LUTG0("~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+~B*A*C*D+B*A*C*D"),
    //.LUTG1("~B*~C*~A*~D+B*~C*~A*~D+~B*C*~A*~D+B*C*~A*~D+~B*~C*A*~D+B*~C*A*~D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011111111),
    .INIT_LUTF1(16'b0101111101011111),
    .INIT_LUTG0(16'b1010000011110000),
    .INIT_LUTG1(16'b0000000001011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg0_b3|t/a/mem_wb/reg2_b3  (
    .a({\t/a/aluin/n12_lutinv ,\t/a/MEM_rd [4]}),
    .c({\t/a/EX_rd [3],\t/a/EX_rs2 [3]}),
    .clk(clock_pad),
    .d({_al_u1984_o,\t/a/EX_rs2 [4]}),
    .e({\t/a/EX_rs2 [3],\t/a/MEM_rd [3]}),
    .mi({\t/a/EX_rd [3],\t/a/MEM_rd [3]}),
    .sr(rst_pad),
    .f({_al_u2010_o,_al_u1970_o}),
    .q({\t/a/MEM_rd [3],\t/a/WB_rd [3]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(~(D*B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b0001001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg0_b4|t/a/id_ex/reg3_b4  (
    .a({\t/a/aluin/n12_lutinv ,\t/a/aluin/sel1_b24/B9 }),
    .b({_al_u1984_o,_al_u2007_o}),
    .c({\t/a/EX_rd [4],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_rs2 [4],\t/a/EX_rs2 [4]}),
    .mi({\t/a/EX_rd [4],\t/a/ID_rs2 [4]}),
    .sr(rst_pad),
    .f({_al_u2000_o,\t/a/EX_B [24]}),
    .q({\t/a/MEM_rd [4],\t/a/EX_rs2 [4]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b0000101001011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg1_b2|t/a/id_ex/reg0_b2  (
    .a({\t/a/alu_B_select [0],_al_u1049_o}),
    .b({open_n32421,_al_u1248_o}),
    .c({\t/a/MEM_aludat [2],_al_u1258_o}),
    .clk(clock_pad),
    .d({\t/a/EX_regdat2 [2],\t/a/reg_writedat [2]}),
    .mi({\t/a/EX_regdat2 [2],open_n32433}),
    .sr(rst_pad),
    .f({_al_u2092_o,\t/a/ID_read_dat2 [2]}),
    .q({\t/a/MEM_regdat2 [2],\t/a/EX_regdat2 [2]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(~C*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg2_b1|t/a/id_ex/reg6_b1  (
    .a({open_n32437,_al_u1747_o}),
    .b({\t/a/EX_op [0],\t/a/ID_op [0]}),
    .c({\t/a/EX_op [2],\t/a/ID_op [1]}),
    .clk(clock_pad),
    .d({\t/a/EX_op [1],\t/a/ID_op [2]}),
    .mi({\t/a/EX_op [1],\t/a/ID_op [1]}),
    .sr(rst_pad),
    .f({_al_u1739_o,\t/a/condition/sel1/B2 }),
    .q({\t/a/MEM_op [1],\t/a/EX_op [1]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*C*D)"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D"),
    //.LUTG0("(A*C*D)"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010000000000000),
    .INIT_LUTF1(16'b0000000001010101),
    .INIT_LUTG0(16'b1010000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg2_b2|t/a/ex_mem/reg2_b0  (
    .a({\t/a/MEM_op [1],\t/a/EX_op [2]}),
    .c({open_n32454,\t/a/EX_op [1]}),
    .clk(clock_pad),
    .d({\t/a/MEM_op [0],\t/a/EX_op [0]}),
    .e({\t/a/MEM_op [2],open_n32456}),
    .mi({\t/a/EX_op [2],\t/a/EX_op [0]}),
    .sr(rst_pad),
    .f({_al_u290_o,_al_u1801_o}),
    .q({\t/a/MEM_op [2],\t/a/MEM_op [0]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*C*~B*A)"),
    //.LUTF1("A*~C*~B*~D+A*C*~B*~D"),
    //.LUTG0("(~1*D*C*~B*A)"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b0000000000100010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg2_b3|t/a/id_ex/reg6_b6  (
    .a({_al_u1739_o,_al_u1739_o}),
    .b({\t/a/EX_op [5],\t/a/EX_op [3]}),
    .c({open_n32472,\t/a/EX_op [4]}),
    .clk(clock_pad),
    .d(\t/a/EX_op [6:5]),
    .e({\t/a/EX_op [3],\t/a/EX_op [6]}),
    .mi({\t/a/EX_op [3],\t/a/ID_op [6]}),
    .sr(rst_pad),
    .f({_al_u1984_o,\t/a/aluin/n10_lutinv }),
    .q({\t/a/MEM_op [3],\t/a/EX_op [6]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*B*A)"),
    //.LUTF1("~C*B*D*~A+C*B*D*~A+~C*B*D*A+C*B*D*A"),
    //.LUTG0("(~1*~D*~C*B*A)"),
    //.LUTG1("C*~B*D*~A+~C*B*D*~A+C*B*D*~A+C*~B*D*A+~C*B*D*A+C*B*D*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b1100110000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg3_b2|t/a/id_ex/reg1_b2  (
    .a({open_n32489,\t/a/aluin/n35_lutinv }),
    .b({\t/a/aluin/n10_lutinv ,\t/a/aluin/n10_lutinv }),
    .c({_al_u1984_o,\t/a/EX_fun3 [0]}),
    .clk(clock_pad),
    .d(\t/a/EX_fun3 [2:1]),
    .e({\t/a/EX_op [4],\t/a/EX_fun3 [2]}),
    .mi({\t/a/EX_fun3 [2],\t/a/ID_fun3 [2]}),
    .sr(rst_pad),
    .f({\t/a/EX_operation [2],_al_u2126_o}),
    .q({\t/a/MEM_fun3 [2],\t/a/EX_fun3 [2]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(~C*~(~D*~A))))"),
    //.LUT1("(B*~(1*~(~C*~(~D*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000110000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b1  (
    .a({\t/a/alu/mux0_b1/B1_0 ,\t/a/alu/mux0_b1/B1_0 }),
    .b({_al_u2586_o,_al_u2586_o}),
    .c({_al_u2587_o,_al_u2587_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n32517,_al_u2128_o}),
    .sr(rst_pad),
    .fx({open_n32521,\t/a/aludat [1]}),
    .q({open_n32522,\t/a/MEM_aludat [1]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b10  (
    .a({_al_u2478_o,_al_u2478_o}),
    .b({_al_u2480_o,_al_u2480_o}),
    .c({_al_u2486_o,_al_u2486_o}),
    .clk(clock_pad),
    .d({_al_u2279_o,_al_u2279_o}),
    .mi({open_n32534,_al_u2161_o}),
    .sr(rst_pad),
    .q({open_n32540,\t/a/MEM_aludat [10]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b11  (
    .a({_al_u2468_o,_al_u2468_o}),
    .b({_al_u2470_o,_al_u2470_o}),
    .c({_al_u2476_o,_al_u2476_o}),
    .clk(clock_pad),
    .d({_al_u2262_o,_al_u2262_o}),
    .mi({open_n32552,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n32556,\t/a/aludat [11]}),
    .q({open_n32557,\t/a/MEM_aludat [11]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b12  (
    .a({_al_u2458_o,_al_u2458_o}),
    .b({_al_u2460_o,_al_u2460_o}),
    .c({_al_u2466_o,_al_u2466_o}),
    .clk(clock_pad),
    .d({_al_u2242_o,_al_u2242_o}),
    .mi({open_n32569,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n32573,\t/a/aludat [12]}),
    .q({open_n32574,\t/a/MEM_aludat [12]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b13  (
    .a({_al_u2448_o,_al_u2448_o}),
    .b({_al_u2450_o,_al_u2450_o}),
    .c({_al_u2456_o,_al_u2456_o}),
    .clk(clock_pad),
    .d({_al_u2219_o,_al_u2219_o}),
    .mi({open_n32586,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n32590,\t/a/aludat [13]}),
    .q({open_n32591,\t/a/MEM_aludat [13]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b14  (
    .a({_al_u2438_o,_al_u2438_o}),
    .b({_al_u2440_o,_al_u2440_o}),
    .c({_al_u2446_o,_al_u2446_o}),
    .clk(clock_pad),
    .d({_al_u2187_o,_al_u2187_o}),
    .mi({open_n32603,_al_u2161_o}),
    .sr(rst_pad),
    .q({open_n32609,\t/a/MEM_aludat [14]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b17  (
    .a({_al_u2405_o,_al_u2405_o}),
    .b({_al_u2406_o,_al_u2406_o}),
    .c({_al_u2412_o,_al_u2412_o}),
    .clk(clock_pad),
    .d({_al_u2413_o,_al_u2413_o}),
    .mi({open_n32621,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32625,\t/a/aludat [17]}),
    .q({open_n32626,\t/a/MEM_aludat [17]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~(0*~A))))"),
    //.LUT1("~(~D*~(C*~(B*~(1*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1111111101110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b18  (
    .a({_al_u2392_o,_al_u2392_o}),
    .b({_al_u2393_o,_al_u2393_o}),
    .c({_al_u2399_o,_al_u2399_o}),
    .clk(clock_pad),
    .d({_al_u2400_o,_al_u2400_o}),
    .mi({open_n32638,_al_u2128_o}),
    .sr(rst_pad),
    .fx({open_n32642,\t/a/aludat [18]}),
    .q({open_n32643,\t/a/MEM_aludat [18]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~(0*~A))))"),
    //.LUT1("~(~D*~(C*~(B*~(1*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1111111101110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b19  (
    .a({_al_u2380_o,_al_u2380_o}),
    .b({_al_u2381_o,_al_u2381_o}),
    .c({_al_u2387_o,_al_u2387_o}),
    .clk(clock_pad),
    .d({_al_u2388_o,_al_u2388_o}),
    .mi({open_n32655,_al_u2128_o}),
    .sr(rst_pad),
    .fx({open_n32659,\t/a/aludat [19]}),
    .q({open_n32660,\t/a/MEM_aludat [19]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(~C*~(~D*~A))))"),
    //.LUT1("(B*~(1*~(~C*~(~D*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000110000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b2  (
    .a({\t/a/alu/mux0_b2/B1_0 ,\t/a/alu/mux0_b2/B1_0 }),
    .b({_al_u2564_o,_al_u2564_o}),
    .c({_al_u2565_o,_al_u2565_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n32672,_al_u2128_o}),
    .sr(rst_pad),
    .fx({open_n32676,\t/a/aludat [2]}),
    .q({open_n32677,\t/a/MEM_aludat [2]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b20  (
    .a({_al_u2368_o,_al_u2368_o}),
    .b({_al_u2369_o,_al_u2369_o}),
    .c({_al_u2375_o,_al_u2375_o}),
    .clk(clock_pad),
    .d({_al_u2376_o,_al_u2376_o}),
    .mi({open_n32689,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32693,\t/a/aludat [20]}),
    .q({open_n32694,\t/a/MEM_aludat [20]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b21  (
    .a({_al_u2355_o,_al_u2355_o}),
    .b({_al_u2356_o,_al_u2356_o}),
    .c({_al_u2362_o,_al_u2362_o}),
    .clk(clock_pad),
    .d({_al_u2363_o,_al_u2363_o}),
    .mi({open_n32706,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32710,\t/a/aludat [21]}),
    .q({open_n32711,\t/a/MEM_aludat [21]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b22  (
    .a({_al_u2342_o,_al_u2342_o}),
    .b({_al_u2343_o,_al_u2343_o}),
    .c({_al_u2349_o,_al_u2349_o}),
    .clk(clock_pad),
    .d({_al_u2350_o,_al_u2350_o}),
    .mi({open_n32723,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32727,\t/a/aludat [22]}),
    .q({open_n32728,\t/a/MEM_aludat [22]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b23  (
    .a({_al_u2329_o,_al_u2329_o}),
    .b({_al_u2330_o,_al_u2330_o}),
    .c({_al_u2336_o,_al_u2336_o}),
    .clk(clock_pad),
    .d({_al_u2337_o,_al_u2337_o}),
    .mi({open_n32740,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32744,\t/a/aludat [23]}),
    .q({open_n32745,\t/a/MEM_aludat [23]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b24  (
    .a({_al_u2310_o,_al_u2310_o}),
    .b({_al_u2317_o,_al_u2317_o}),
    .c({_al_u2323_o,_al_u2323_o}),
    .clk(clock_pad),
    .d({_al_u2324_o,_al_u2324_o}),
    .mi({open_n32757,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32761,\t/a/aludat [24]}),
    .q({open_n32762,\t/a/MEM_aludat [24]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b25  (
    .a({_al_u2293_o,_al_u2293_o}),
    .b({_al_u2301_o,_al_u2301_o}),
    .c({_al_u2307_o,_al_u2307_o}),
    .clk(clock_pad),
    .d({_al_u2308_o,_al_u2308_o}),
    .mi({open_n32774,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32778,\t/a/aludat [25]}),
    .q({open_n32779,\t/a/MEM_aludat [25]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b26  (
    .a({_al_u2276_o,_al_u2276_o}),
    .b({_al_u2284_o,_al_u2284_o}),
    .c({_al_u2290_o,_al_u2290_o}),
    .clk(clock_pad),
    .d({_al_u2291_o,_al_u2291_o}),
    .mi({open_n32791,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32795,\t/a/aludat [26]}),
    .q({open_n32796,\t/a/MEM_aludat [26]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b27  (
    .a({_al_u2259_o,_al_u2259_o}),
    .b({_al_u2267_o,_al_u2267_o}),
    .c({_al_u2273_o,_al_u2273_o}),
    .clk(clock_pad),
    .d({_al_u2274_o,_al_u2274_o}),
    .mi({open_n32808,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32812,\t/a/aludat [27]}),
    .q({open_n32813,\t/a/MEM_aludat [27]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b28  (
    .a({_al_u2236_o,_al_u2236_o}),
    .b({_al_u2250_o,_al_u2250_o}),
    .c({_al_u2256_o,_al_u2256_o}),
    .clk(clock_pad),
    .d({_al_u2257_o,_al_u2257_o}),
    .mi({open_n32825,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32829,\t/a/aludat [28]}),
    .q({open_n32830,\t/a/MEM_aludat [28]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b29  (
    .a({_al_u2212_o,_al_u2212_o}),
    .b({_al_u2227_o,_al_u2227_o}),
    .c({_al_u2233_o,_al_u2233_o}),
    .clk(clock_pad),
    .d({_al_u2234_o,_al_u2234_o}),
    .mi({open_n32842,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32846,\t/a/aludat [29]}),
    .q({open_n32847,\t/a/MEM_aludat [29]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(~C*~(~D*~A))))"),
    //.LUT1("(B*~(1*~(~C*~(~D*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000110000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b3  (
    .a({\t/a/alu/mux0_b3/B1_0 ,\t/a/alu/mux0_b3/B1_0 }),
    .b({_al_u2555_o,_al_u2555_o}),
    .c({_al_u2556_o,_al_u2556_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n32859,_al_u2128_o}),
    .sr(rst_pad),
    .q({open_n32865,\t/a/MEM_aludat [3]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b30  (
    .a({_al_u2172_o,_al_u2172_o}),
    .b({_al_u2203_o,_al_u2203_o}),
    .c({_al_u2209_o,_al_u2209_o}),
    .clk(clock_pad),
    .d({_al_u2210_o,_al_u2210_o}),
    .mi({open_n32877,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32881,\t/a/aludat [30]}),
    .q({open_n32882,\t/a/MEM_aludat [30]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b31  (
    .a({_al_u2130_o,_al_u2130_o}),
    .b({_al_u2163_o,_al_u2163_o}),
    .c({_al_u2168_o,_al_u2168_o}),
    .clk(clock_pad),
    .d({_al_u2170_o,_al_u2170_o}),
    .mi({open_n32894,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n32898,\t/a/aludat [31]}),
    .q({open_n32899,\t/a/MEM_aludat [31]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(~C*~(~D*~A))))"),
    //.LUT1("(A*~(1*~(~C*~(~D*~B))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000101000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b5  (
    .a({_al_u2535_o,\t/a/alu/mux0_b5/B1_0 }),
    .b({\t/a/alu/mux0_b5/B1_0 ,_al_u2535_o}),
    .c({_al_u2536_o,_al_u2536_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n32911,_al_u2128_o}),
    .sr(rst_pad),
    .q({open_n32917,\t/a/MEM_aludat [5]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(~C*~(~D*~A))))"),
    //.LUT1("(B*~(1*~(~C*~(~D*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000110000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b6  (
    .a({\t/a/alu/mux0_b6/B1_0 ,\t/a/alu/mux0_b6/B1_0 }),
    .b({_al_u2525_o,_al_u2525_o}),
    .c({_al_u2526_o,_al_u2526_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n32929,_al_u2128_o}),
    .sr(rst_pad),
    .q({open_n32935,\t/a/MEM_aludat [6]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*D)))"),
    //.LUT1("(~C*B*~(A*~(1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000110000000100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b7  (
    .a({_al_u2508_o,_al_u2508_o}),
    .b({_al_u2510_o,_al_u2510_o}),
    .c({_al_u2516_o,_al_u2516_o}),
    .clk(clock_pad),
    .d({\t/a/alu/n260_lutinv ,\t/a/alu/n260_lutinv }),
    .mi({open_n32947,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n32951,\t/a/aludat [7]}),
    .q({open_n32952,\t/a/MEM_aludat [7]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b8  (
    .a({_al_u2498_o,_al_u2498_o}),
    .b({_al_u2500_o,_al_u2500_o}),
    .c({_al_u2506_o,_al_u2506_o}),
    .clk(clock_pad),
    .d({_al_u2312_o,_al_u2312_o}),
    .mi({open_n32964,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n32968,\t/a/aludat [8]}),
    .q({open_n32969,\t/a/MEM_aludat [8]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b9  (
    .a({_al_u2488_o,_al_u2488_o}),
    .b({_al_u2490_o,_al_u2490_o}),
    .c({_al_u2496_o,_al_u2496_o}),
    .clk(clock_pad),
    .d({_al_u2296_o,_al_u2296_o}),
    .mi({open_n32981,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n32985,\t/a/aludat [9]}),
    .q({open_n32986,\t/a/MEM_aludat [9]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~C*~A*~D+B*~C*~A*~D+~B*C*~A*~D+B*C*~A*~D+~B*~C*A*~D+~B*C*A*~D+B*~C*~A*D+B*C*~A*D"),
    //.LUTF1("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+A*~C*B*~D+A*C*B*~D+A*~C*B*D+A*C*B*D"),
    //.LUTG0("0"),
    //.LUTG1("A*~C*B*~D+A*C*B*~D+A*~C*B*D+A*C*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010001110111),
    .INIT_LUTF1(16'b1000100010111011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b0|t/a/ex_mem/reg1_b0  (
    .a({\t/a/reg_writedat [0],\t/a/MEM_aludat [0]}),
    .b({_al_u1049_o,\t/a/alu_B_select [0]}),
    .clk(clock_pad),
    .d({_al_u1720_o,\t/a/EX_regdat2 [0]}),
    .e({_al_u1710_o,\t/a/alu_B_select [1]}),
    .mi({open_n32991,\t/a/EX_regdat2 [0]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [0],_al_u2075_o}),
    .q({\t/a/EX_regdat2 [0],\t/a/MEM_regdat2 [0]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1100110100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b10|t/a/ex_mem/reg1_b10  (
    .a({_al_u1689_o,\t/a/alu_B_select [0]}),
    .b({_al_u1049_o,\t/a/alu_B_select [1]}),
    .c({_al_u1699_o,\t/a/MEM_aludat [10]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [10],\t/a/EX_regdat2 [10]}),
    .mi({open_n33017,\t/a/EX_regdat2 [10]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [10],_al_u2069_o}),
    .q({\t/a/EX_regdat2 [10],\t/a/MEM_regdat2 [10]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~D*~A)*~(C)*~(B)+(~D*~A)*C*~(B)+~((~D*~A))*C*B+(~D*~A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1100000011010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b11|t/a/ex_mem/reg1_b11  (
    .a({_al_u1668_o,\t/a/alu_B_select [0]}),
    .b({_al_u1049_o,\t/a/alu_B_select [1]}),
    .c({\t/a/reg_writedat [11],\t/a/MEM_aludat [11]}),
    .clk(clock_pad),
    .d({_al_u1678_o,\t/a/EX_regdat2 [11]}),
    .mi({open_n33032,\t/a/EX_regdat2 [11]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [11],_al_u2066_o}),
    .q({\t/a/EX_regdat2 [11],\t/a/MEM_regdat2 [11]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~C*~A*~D+B*~C*~A*~D+~B*C*~A*~D+B*C*~A*~D+~B*~C*A*~D+~B*C*A*~D+B*~C*~A*D+B*C*~A*D"),
    //.LUTF1("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D+C*~B*~A*D+C*B*~A*D+C*~B*A*D+C*B*A*D"),
    //.LUTG0("0"),
    //.LUTG1("C*~B*~A*D+C*B*~A*D+C*~B*A*D+C*B*A*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010001110111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b12|t/a/ex_mem/reg1_b12  (
    .a({open_n33036,\t/a/MEM_aludat [12]}),
    .b({_al_u1647_o,\t/a/alu_B_select [0]}),
    .c({\t/a/reg_writedat [12],open_n33037}),
    .clk(clock_pad),
    .d({_al_u1049_o,\t/a/EX_regdat2 [12]}),
    .e({_al_u1657_o,\t/a/alu_B_select [1]}),
    .mi({open_n33040,\t/a/EX_regdat2 [12]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [12],_al_u2063_o}),
    .q({\t/a/EX_regdat2 [12],\t/a/MEM_regdat2 [12]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D"),
    //.LUTG0("~A*~B*~C*~D+~A*~B*C*~D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000110011),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000000000010001),
    .INIT_LUTG1(16'b1111000011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b13|t/a/ex_mem/reg1_b13  (
    .a({open_n33055,\t/a/alu_B_select [0]}),
    .b({_al_u1626_o,\t/a/alu_B_select [1]}),
    .c({_al_u1049_o,open_n33056}),
    .clk(clock_pad),
    .d({_al_u1636_o,\t/a/EX_regdat2 [13]}),
    .e({\t/a/reg_writedat [13],\t/a/MEM_aludat [13]}),
    .mi({open_n33059,\t/a/EX_regdat2 [13]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [13],_al_u2060_o}),
    .q({\t/a/EX_regdat2 [13],\t/a/MEM_regdat2 [13]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1100110100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b14|t/a/ex_mem/reg1_b14  (
    .a({_al_u1605_o,\t/a/alu_B_select [0]}),
    .b({_al_u1049_o,\t/a/alu_B_select [1]}),
    .c({_al_u1615_o,\t/a/MEM_aludat [14]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [14],\t/a/EX_regdat2 [14]}),
    .mi({open_n33085,\t/a/EX_regdat2 [14]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [14],_al_u2057_o}),
    .q({\t/a/EX_regdat2 [14],\t/a/MEM_regdat2 [14]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1100110100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b15|t/a/ex_mem/reg1_b15  (
    .a({_al_u1584_o,\t/a/alu_B_select [0]}),
    .b({_al_u1049_o,\t/a/alu_B_select [1]}),
    .c({_al_u1594_o,\t/a/MEM_aludat [15]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [15],\t/a/EX_regdat2 [15]}),
    .mi({open_n33100,\t/a/EX_regdat2 [15]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [15],_al_u2054_o}),
    .q({\t/a/EX_regdat2 [15],\t/a/MEM_regdat2 [15]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~B*~C*~D+~A*~B*C*~D"),
    //.LUTG1("~A*B*C*~D+A*B*C*~D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000110011),
    .INIT_LUTF1(16'b1100000011001111),
    .INIT_LUTG0(16'b0000000000010001),
    .INIT_LUTG1(16'b1100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b16|t/a/ex_mem/reg1_b16  (
    .a({open_n33104,\t/a/alu_B_select [0]}),
    .b({\t/a/reg_writedat [16],\t/a/alu_B_select [1]}),
    .c({_al_u1049_o,open_n33105}),
    .clk(clock_pad),
    .d({_al_u1563_o,\t/a/EX_regdat2 [16]}),
    .e({_al_u1573_o,\t/a/MEM_aludat [16]}),
    .mi({open_n33108,\t/a/EX_regdat2 [16]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [16],_al_u2051_o}),
    .q({\t/a/EX_regdat2 [16],\t/a/MEM_regdat2 [16]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+A*~C*~B*D+A*C*~B*D"),
    //.LUTF1("~D*~A*~C*~B+D*~A*~C*~B+~D*A*~C*~B+D*A*~C*~B+D*~A*~C*B+D*A*~C*B+D*~A*C*B+D*A*C*B"),
    //.LUTG0("0"),
    //.LUTG1("D*~A*~C*B+D*A*~C*B+D*~A*C*B+D*A*C*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001001110111),
    .INIT_LUTF1(16'b1100111100000011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1100110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b17|t/a/ex_mem/reg1_b17  (
    .a({open_n33123,\t/a/alu_B_select [0]}),
    .b({_al_u1049_o,\t/a/MEM_aludat [17]}),
    .c({_al_u1552_o,open_n33124}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [17],\t/a/EX_regdat2 [17]}),
    .e({_al_u1542_o,\t/a/alu_B_select [1]}),
    .mi({open_n33127,\t/a/EX_regdat2 [17]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [17],_al_u2048_o}),
    .q({\t/a/EX_regdat2 [17],\t/a/MEM_regdat2 [17]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b18|t/a/ex_mem/reg1_b18  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1521_o,\t/a/alu_B_select [1]}),
    .c({_al_u1531_o,\t/a/MEM_aludat [18]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [18],\t/a/EX_regdat2 [18]}),
    .mi({open_n33153,\t/a/EX_regdat2 [18]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [18],_al_u2045_o}),
    .q({\t/a/EX_regdat2 [18],\t/a/MEM_regdat2 [18]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b19|t/a/ex_mem/reg1_b19  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1500_o,\t/a/alu_B_select [1]}),
    .c({_al_u1510_o,\t/a/MEM_aludat [19]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [19],\t/a/EX_regdat2 [19]}),
    .mi({open_n33168,\t/a/EX_regdat2 [19]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [19],_al_u2042_o}),
    .q({\t/a/EX_regdat2 [19],\t/a/MEM_regdat2 [19]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*~C*~D+B*~A*~C*~D+~B*~A*C*~D+B*~A*C*~D"),
    //.LUTF1("~D*~A*~C*~B+D*~A*~C*~B+~D*A*~C*~B+D*A*~C*~B+D*~A*~C*B+D*A*~C*B+D*~A*C*B+D*A*C*B"),
    //.LUTG0("~B*~A*~C*~D+B*~A*~C*~D+~B*~A*~C*D+B*~A*~C*D"),
    //.LUTG1("D*~A*~C*B+D*A*~C*B+D*~A*C*B+D*A*C*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000001010101),
    .INIT_LUTF1(16'b1100111100000011),
    .INIT_LUTG0(16'b0000010100000101),
    .INIT_LUTG1(16'b1100110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b1|t/a/ex_mem/reg1_b1  (
    .a({open_n33172,\t/a/alu_B_select [1]}),
    .b({_al_u1049_o,open_n33173}),
    .c({_al_u1489_o,\t/a/MEM_aludat [1]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [1],\t/a/EX_regdat2 [1]}),
    .e({_al_u1479_o,\t/a/alu_B_select [0]}),
    .mi({open_n33176,\t/a/EX_regdat2 [1]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [1],_al_u2072_o}),
    .q({\t/a/EX_regdat2 [1],\t/a/MEM_regdat2 [1]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~C*~A*~D+B*~C*~A*~D+~B*C*~A*~D+B*C*~A*~D+~B*~C*A*~D+~B*C*A*~D+B*~C*~A*D+B*C*~A*D"),
    //.LUTF1("((~A*~B)*~(D)*~(C)+(~A*~B)*D*~(C)+~((~A*~B))*D*C+(~A*~B)*D*C)"),
    //.LUTG0("0"),
    //.LUTG1("((~A*~B)*~(D)*~(C)+(~A*~B)*D*~(C)+~((~A*~B))*D*C+(~A*~B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010001110111),
    .INIT_LUTF1(16'b1111000100000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b20|t/a/ex_mem/reg1_b20  (
    .a({_al_u1468_o,\t/a/MEM_aludat [20]}),
    .b({_al_u1458_o,\t/a/alu_B_select [0]}),
    .c({_al_u1049_o,open_n33191}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [20],\t/a/EX_regdat2 [20]}),
    .e({open_n33193,\t/a/alu_B_select [1]}),
    .mi({open_n33195,\t/a/EX_regdat2 [20]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [20],_al_u2039_o}),
    .q({\t/a/EX_regdat2 [20],\t/a/MEM_regdat2 [20]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*~B*~C*D+A*B*~C*D"),
    //.LUTF1("~A*~C*~D*~B+~A*C*~D*~B+~A*C*D*~B+A*C*D*~B+~A*~C*~D*B+~A*C*~D*B+~A*C*D*B+A*C*D*B"),
    //.LUTG0("0"),
    //.LUTG1("~A*C*D*~B+A*C*D*~B+~A*C*D*B+A*C*D*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101001011111),
    .INIT_LUTF1(16'b1111000001010101),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b21|t/a/ex_mem/reg1_b21  (
    .a({_al_u1447_o,\t/a/alu_B_select [0]}),
    .c({\t/a/reg_writedat [21],\t/a/MEM_aludat [21]}),
    .clk(clock_pad),
    .d({_al_u1049_o,\t/a/EX_regdat2 [21]}),
    .e({_al_u1437_o,\t/a/alu_B_select [1]}),
    .mi({open_n33214,\t/a/EX_regdat2 [21]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [21],_al_u2036_o}),
    .q({\t/a/EX_regdat2 [21],\t/a/MEM_regdat2 [21]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~D*~B)*~(C)*~(A)+(~D*~B)*C*~(A)+~((~D*~B))*C*A+(~D*~B)*C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010000010110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b22|t/a/ex_mem/reg1_b22  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1416_o,\t/a/alu_B_select [1]}),
    .c({\t/a/reg_writedat [22],\t/a/MEM_aludat [22]}),
    .clk(clock_pad),
    .d({_al_u1426_o,\t/a/EX_regdat2 [22]}),
    .mi({open_n33240,\t/a/EX_regdat2 [22]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [22],_al_u2033_o}),
    .q({\t/a/EX_regdat2 [22],\t/a/MEM_regdat2 [22]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~D)*~(B)*~(A)+(~C*~D)*B*~(A)+~((~C*~D))*B*A+(~C*~D)*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1000100010001101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b23|t/a/ex_mem/reg1_b23  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({\t/a/reg_writedat [23],\t/a/alu_B_select [1]}),
    .c({_al_u1405_o,\t/a/MEM_aludat [23]}),
    .clk(clock_pad),
    .d({_al_u1395_o,\t/a/EX_regdat2 [23]}),
    .mi({open_n33255,\t/a/EX_regdat2 [23]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [23],_al_u2030_o}),
    .q({\t/a/EX_regdat2 [23],\t/a/MEM_regdat2 [23]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*~B*~C*D+A*B*~C*D"),
    //.LUTF1("~A*~C*~D*~B+A*~C*~D*~B+~A*~C*D*~B+A*~C*D*~B+A*~C*~D*B+A*C*~D*B+A*~C*D*B+A*C*D*B"),
    //.LUTG0("0"),
    //.LUTG1("A*~C*~D*B+A*C*~D*B+A*~C*D*B+A*C*D*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101001011111),
    .INIT_LUTF1(16'b1000101110001011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1000100010001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b24|t/a/ex_mem/reg1_b24  (
    .a({\t/a/reg_writedat [24],\t/a/alu_B_select [0]}),
    .b({_al_u1049_o,open_n33259}),
    .c({_al_u1374_o,\t/a/MEM_aludat [24]}),
    .clk(clock_pad),
    .d({open_n33261,\t/a/EX_regdat2 [24]}),
    .e({_al_u1384_o,\t/a/alu_B_select [1]}),
    .mi({open_n33263,\t/a/EX_regdat2 [24]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [24],_al_u2027_o}),
    .q({\t/a/EX_regdat2 [24],\t/a/MEM_regdat2 [24]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*~B*~C*D+A*B*~C*D"),
    //.LUTF1("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D+C*~B*~A*D+C*B*~A*D+C*~B*A*D+C*B*A*D"),
    //.LUTG0("0"),
    //.LUTG1("C*~B*~A*D+C*B*~A*D+C*~B*A*D+C*B*A*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101001011111),
    .INIT_LUTF1(16'b1111000000110011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b25|t/a/ex_mem/reg1_b25  (
    .a({open_n33278,\t/a/alu_B_select [0]}),
    .b({_al_u1353_o,open_n33279}),
    .c({\t/a/reg_writedat [25],\t/a/MEM_aludat [25]}),
    .clk(clock_pad),
    .d({_al_u1049_o,\t/a/EX_regdat2 [25]}),
    .e({_al_u1363_o,\t/a/alu_B_select [1]}),
    .mi({open_n33282,\t/a/EX_regdat2 [25]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [25],_al_u2024_o}),
    .q({\t/a/EX_regdat2 [25],\t/a/MEM_regdat2 [25]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1100110100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b26|t/a/ex_mem/reg1_b26  (
    .a({_al_u1332_o,\t/a/alu_B_select [0]}),
    .b({_al_u1049_o,\t/a/alu_B_select [1]}),
    .c({_al_u1342_o,\t/a/MEM_aludat [26]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [26],\t/a/EX_regdat2 [26]}),
    .mi({open_n33308,\t/a/EX_regdat2 [26]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [26],_al_u2021_o}),
    .q({\t/a/EX_regdat2 [26],\t/a/MEM_regdat2 [26]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~D)*~(A)*~(B)+(~C*~D)*A*~(B)+~((~C*~D))*A*B+(~C*~D)*A*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1000100010001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b27|t/a/ex_mem/reg1_b27  (
    .a({\t/a/reg_writedat [27],\t/a/alu_B_select [0]}),
    .b({_al_u1049_o,\t/a/alu_B_select [1]}),
    .c({_al_u1321_o,\t/a/MEM_aludat [27]}),
    .clk(clock_pad),
    .d({_al_u1311_o,\t/a/EX_regdat2 [27]}),
    .mi({open_n33323,\t/a/EX_regdat2 [27]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [27],_al_u2018_o}),
    .q({\t/a/EX_regdat2 [27],\t/a/MEM_regdat2 [27]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*B*~D+~A*C*B*~D+A*~C*~B*D+A*C*~B*D"),
    //.LUTF1("~C*~A*~B*~D+C*~A*~B*~D+~C*A*~B*~D+C*A*~B*~D+C*~A*B*~D+C*A*B*~D+C*~A*B*D+C*A*B*D"),
    //.LUTG0("0"),
    //.LUTG1("C*~A*B*~D+C*A*B*~D+C*~A*B*D+C*A*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001001110111),
    .INIT_LUTF1(16'b1100000011110011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b28|t/a/ex_mem/reg1_b28  (
    .a({open_n33327,\t/a/alu_B_select [0]}),
    .b({_al_u1049_o,\t/a/MEM_aludat [28]}),
    .c({\t/a/reg_writedat [28],open_n33328}),
    .clk(clock_pad),
    .d({_al_u1300_o,\t/a/EX_regdat2 [28]}),
    .e({_al_u1290_o,\t/a/alu_B_select [1]}),
    .mi({open_n33331,\t/a/EX_regdat2 [28]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [28],_al_u2015_o}),
    .q({\t/a/EX_regdat2 [28],\t/a/MEM_regdat2 [28]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*~B*~C*A+D*~B*~C*A"),
    //.LUTG0("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*~A*D+C*~B*~A*D"),
    //.LUTG1("D*~B*~C*~A+D*B*~C*~A+D*~B*C*~A+D*B*C*~A+D*~B*~C*A+D*B*~C*A+D*~B*C*A+D*B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000110011),
    .INIT_LUTF1(16'b0000001100000011),
    .INIT_LUTG0(16'b0001000100010001),
    .INIT_LUTG1(16'b1111111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b29|t/a/ex_mem/reg1_b29  (
    .a({open_n33346,\t/a/MEM_aludat [29]}),
    .b({_al_u1269_o,\t/a/alu_B_select [1]}),
    .c({_al_u1279_o,open_n33347}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [29],\t/a/EX_regdat2 [29]}),
    .e({_al_u1049_o,\t/a/alu_B_select [0]}),
    .mi({open_n33350,\t/a/EX_regdat2 [29]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [29],_al_u2012_o}),
    .q({\t/a/EX_regdat2 [29],\t/a/MEM_regdat2 [29]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b30|t/a/ex_mem/reg1_b30  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1227_o,\t/a/alu_B_select [1]}),
    .c({_al_u1237_o,\t/a/MEM_aludat [30]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [30],\t/a/EX_regdat2 [30]}),
    .mi({open_n33376,\t/a/EX_regdat2 [30]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [30],_al_u2005_o}),
    .q({\t/a/EX_regdat2 [30],\t/a/MEM_regdat2 [30]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+~B*~A*C*~D+~B*A*C*~D+B*~A*~C*D+B*A*~C*D"),
    //.LUTF1("~B*~A*~C*~D+~B*A*~C*~D+~B*~A*~C*D+~B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    //.LUTG0("0"),
    //.LUTG1("~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000110000111111),
    .INIT_LUTF1(16'b1111001100000011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b31|t/a/ex_mem/reg1_b31  (
    .b({_al_u1216_o,\t/a/alu_B_select [0]}),
    .c({_al_u1049_o,\t/a/MEM_aludat [31]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [31],\t/a/EX_regdat2 [31]}),
    .e({_al_u1206_o,\t/a/alu_B_select [1]}),
    .mi({open_n33384,\t/a/EX_regdat2 [31]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [31],_al_u2002_o}),
    .q({\t/a/EX_regdat2 [31],\t/a/MEM_regdat2 [31]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b3|t/a/ex_mem/reg1_b3  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1185_o,\t/a/alu_B_select [1]}),
    .c({_al_u1195_o,\t/a/MEM_aludat [3]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [3],\t/a/EX_regdat2 [3]}),
    .mi({open_n33410,\t/a/EX_regdat2 [3]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [3],_al_u2009_o}),
    .q({\t/a/EX_regdat2 [3],\t/a/MEM_regdat2 [3]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    //.LUTF1("~B*~A*~C*~D+B*~A*~C*~D+~B*A*~C*~D+B*A*~C*~D+B*~A*~C*D+B*A*~C*D+B*~A*C*D+B*A*C*D"),
    //.LUTG0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTG1("B*~A*~C*D+B*A*~C*D+B*~A*C*D+B*A*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000110011),
    .INIT_LUTF1(16'b1100110000001111),
    .INIT_LUTG0(16'b0000001100000011),
    .INIT_LUTG1(16'b1100110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b4|t/a/ex_mem/reg1_b4  (
    .b({\t/a/reg_writedat [4],\t/a/alu_B_select [1]}),
    .c({_al_u1174_o,\t/a/MEM_aludat [4]}),
    .clk(clock_pad),
    .d({_al_u1049_o,\t/a/EX_regdat2 [4]}),
    .e({_al_u1164_o,\t/a/alu_B_select [0]}),
    .mi({open_n33418,\t/a/EX_regdat2 [4]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [4],_al_u1999_o}),
    .q({\t/a/EX_regdat2 [4],\t/a/MEM_regdat2 [4]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b5|t/a/ex_mem/reg1_b5  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1143_o,\t/a/alu_B_select [1]}),
    .c({_al_u1153_o,\t/a/MEM_aludat [5]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [5],\t/a/EX_regdat2 [5]}),
    .mi({open_n33444,\t/a/EX_regdat2 [5]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [5],_al_u1996_o}),
    .q({\t/a/EX_regdat2 [5],\t/a/MEM_regdat2 [5]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1100110100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b6|t/a/ex_mem/reg1_b6  (
    .a({_al_u1122_o,\t/a/alu_B_select [0]}),
    .b({_al_u1049_o,\t/a/alu_B_select [1]}),
    .c({_al_u1132_o,\t/a/MEM_aludat [6]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [6],\t/a/EX_regdat2 [6]}),
    .mi({open_n33459,\t/a/EX_regdat2 [6]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [6],_al_u1993_o}),
    .q({\t/a/EX_regdat2 [6],\t/a/MEM_regdat2 [6]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    //.LUTF1("~C*~A*~B*~D+C*~A*~B*~D+~C*A*~B*~D+C*A*~B*~D+C*~A*B*~D+C*A*B*~D+C*~A*B*D+C*A*B*D"),
    //.LUTG0("~A*~B*~C*~D+~A*~B*C*~D"),
    //.LUTG1("C*~A*B*~D+C*A*B*~D+C*~A*B*D+C*A*B*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000110011),
    .INIT_LUTF1(16'b1100000011110011),
    .INIT_LUTG0(16'b0000000000010001),
    .INIT_LUTG1(16'b1100000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b7|t/a/ex_mem/reg1_b7  (
    .a({open_n33463,\t/a/alu_B_select [0]}),
    .b({_al_u1049_o,\t/a/alu_B_select [1]}),
    .c({\t/a/reg_writedat [7],open_n33464}),
    .clk(clock_pad),
    .d({_al_u1111_o,\t/a/EX_regdat2 [7]}),
    .e({_al_u1101_o,\t/a/MEM_aludat [7]}),
    .mi({open_n33467,\t/a/EX_regdat2 [7]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [7],_al_u1990_o}),
    .q({\t/a/EX_regdat2 [7],\t/a/MEM_regdat2 [7]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*~B*~C*D+A*~B*C*D"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*~B*~C*~D+~A*~B*C*~D"),
    //.LUTG1("~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000110011),
    .INIT_LUTF1(16'b1111010100000101),
    .INIT_LUTG0(16'b0000000000010001),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b8|t/a/ex_mem/reg1_b8  (
    .a({_al_u1090_o,\t/a/alu_B_select [0]}),
    .b({open_n33482,\t/a/alu_B_select [1]}),
    .c({_al_u1049_o,open_n33483}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [8],\t/a/EX_regdat2 [8]}),
    .e({_al_u1080_o,\t/a/MEM_aludat [8]}),
    .mi({open_n33486,\t/a/EX_regdat2 [8]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [8],_al_u1987_o}),
    .q({\t/a/EX_regdat2 [8],\t/a/MEM_regdat2 [8]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~D*~B)*~(C)*~(A)+(~D*~B)*C*~(A)+~((~D*~B))*C*A+(~D*~B)*C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010000010110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b9|t/a/ex_mem/reg1_b9  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1059_o,\t/a/alu_B_select [1]}),
    .c({\t/a/reg_writedat [9],\t/a/MEM_aludat [9]}),
    .clk(clock_pad),
    .d({_al_u1069_o,\t/a/EX_regdat2 [9]}),
    .mi({open_n33512,\t/a/EX_regdat2 [9]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [9],_al_u1979_o}),
    .q({\t/a/EX_regdat2 [9],\t/a/MEM_regdat2 [9]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*(C@(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTF1("(~0*~D*(C@(B*A)))"),
    //.LUTG0("(1*(C@(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTG1("(~1*~D*(C@(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000001111000),
    .INIT_LUTG0(16'b0011110001011010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg1_b0|t/a/id_ex/reg1_b1  (
    .a({_al_u2777_o,\t/a/condition/n9 }),
    .b({_al_u2790_o,\t/a/condition/n10 }),
    .c({\t/a/ID_fun3 [0],\t/a/ID_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/ID_fun3 [1],\t/a/ID_fun3 [1]}),
    .e({\t/a/ID_fun3 [2],\t/a/ID_fun3 [2]}),
    .mi({\t/a/ID_fun3 [0],\t/a/ID_fun3 [1]}),
    .sr(rst_pad),
    .f({_al_u2791_o,_al_u2766_o}),
    .q({\t/a/EX_fun3 [0],\t/a/EX_fun3 [1]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*C)*~(0*A))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~B*~(D*C)*~(1*A))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b1111101010101010),
    .INIT_LUTG0(16'b0000000100010001),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg3_b2|t/a/ex_mem/reg0_b2  (
    .a({\t/a/aluin/sel1_b22/B9 ,\t/a/aluin/n12_lutinv }),
    .b({open_n33532,_al_u1802_o}),
    .c({_al_u1803_o,_al_u1984_o}),
    .clk(clock_pad),
    .d({\t/a/EX_rs2 [2],\t/a/EX_rs2 [2]}),
    .e({_al_u2007_o,\t/a/EX_rd [2]}),
    .mi({\t/a/ID_rs2$2$_placeOpt_7 ,\t/a/EX_rd [2]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [22],_al_u2093_o}),
    .q({\t/a/EX_rs2 [2],\t/a/MEM_rd [2]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("((B@D)*(C@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0001001001001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg5_b0|t/a/if_id/reg2_b0  (
    .a({_al_u2111_o,\t/a/if_id/n9 }),
    .b({\t/a/ID_rd [0],\t/busarbitration/n3_placeOpt_5 }),
    .c({\t/a/ID_rd [4],\t/busarbitration/instruction [7]}),
    .clk(clock_pad),
    .d({_al_u2119_o,i_data[7]}),
    .mi({\t/a/ID_rd [0],open_n33560}),
    .sr(rst_pad),
    .f({_al_u2806_o,open_n33561}),
    .q({\t/a/EX_rd [0],\t/a/ID_rd [0]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1010000010100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg5_b3|t/a/if_id/reg2_b3  (
    .a({_al_u2113_o,\t/a/if_id/n9 }),
    .b({open_n33565,\t/busarbitration/n3_placeOpt_5 }),
    .c({\t/a/ID_rd [3],\t/busarbitration/instruction [10]}),
    .clk(clock_pad),
    .d({open_n33567,i_data[10]}),
    .mi({\t/a/ID_rd [3],open_n33578}),
    .sr(rst_pad),
    .f({_al_u2799_o,open_n33579}),
    .q({\t/a/EX_rd [3],\t/a/ID_rd [3]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~B*C*~A+D*~B*C*~A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTF1("C*B*~A*~D+C*B*A*~D+~C*B*~A*D+~C*B*A*D"),
    //.LUTG0("0"),
    //.LUTG1("C*~B*~A*~D+C*~B*A*~D+~C*~B*~A*D+~C*~B*A*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011100010111000),
    .INIT_LUTF1(16'b0000110011000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000001100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg5_b4|t/a/if_id/reg2_b4  (
    .a({open_n33583,i_data[11]}),
    .b({_al_u1960_o,\t/busarbitration/n3_placeOpt_5 }),
    .c({_al_u1956_o,\t/busarbitration/instruction [11]}),
    .clk(clock_pad),
    .d({\t/a/ID_rd [4],open_n33585}),
    .e({\t/a/ID_rd [2],\t/a/if_id/n9 }),
    .mi({\t/a/ID_rd [4],open_n33587}),
    .sr(rst_pad),
    .f({_al_u2793_o,open_n33599}),
    .q({\t/a/EX_rd [4],\t/a/ID_rd [4]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~D*~C*A*~B+D*~C*A*~B+~D*C*~A*B+D*C*~A*B+~D*~C*A*B+D*~C*A*B+~D*C*A*B+D*C*A*B"),
    //.LUTF1("0"),
    //.LUTG0("0"),
    //.LUTG1("~C*B*D*~A+~C*B*D*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100101011001010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg6_b0|t/a/if_id/reg6_b0  (
    .a({open_n33603,\t/busarbitration/instruction [0]}),
    .b({\t/a/ID_op [1],i_data[0]}),
    .c({\t/a/ID_op [2],\t/busarbitration/n3_placeOpt_2 }),
    .clk(clock_pad),
    .d({\t/a/ID_op [0],open_n33605}),
    .e({_al_u2803_o,\t/a/if_id/n9 }),
    .mi({\t/a/ID_op [0],open_n33607}),
    .sr(rst_pad),
    .f({\t/a/n0_lutinv ,open_n33619}),
    .q({\t/a/EX_op [0],\t/a/ID_op [0]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~C*~B*~D+A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D"),
    //.LUTF1("0"),
    //.LUTG0("0"),
    //.LUTG1("~A*~D*C*B+~A*D*C*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100110011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0100000001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg6_b2|t/a/if_id/reg6_b2  (
    .a({\t/a/ID_op [2],open_n33623}),
    .b({_al_u1747_o,\t/instruction$2$_neg_lutinv }),
    .c({\t/a/ID_op [0],open_n33624}),
    .clk(clock_pad),
    .e({\t/a/ID_op [1],\t/a/if_id/n9 }),
    .mi({\t/a/ID_op [2],open_n33629}),
    .sr(rst_pad),
    .f({\t/a/condition/n1_lutinv ,open_n33641}),
    .q({\t/a/EX_op [2],\t/a/ID_op [2]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg6_b3|t/a/if_id/reg6_b6  (
    .a({\t/a/ID_op [3],\t/a/if_id/n9 }),
    .b({\t/a/ID_op [4],\t/busarbitration/n3_placeOpt_2 }),
    .c({\t/a/ID_op [5],\t/busarbitration/instruction [6]}),
    .clk(clock_pad),
    .d({\t/a/ID_op [6],i_data[6]}),
    .mi({\t/a/ID_op [3],open_n33656}),
    .sr(rst_pad),
    .f({_al_u2803_o,open_n33657}),
    .q({\t/a/EX_op [3],\t/a/ID_op [6]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(C*D*~A*~B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0001000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg6_b4|t/a/if_id/reg6_b5  (
    .a({\t/a/ID_op [4],\t/a/if_id/n9 }),
    .b({\t/a/ID_op [3],\t/busarbitration/n3_placeOpt_2 }),
    .c({\t/a/ID_op [6],\t/busarbitration/instruction [5]}),
    .clk(clock_pad),
    .d({\t/a/ID_op [5],i_data[5]}),
    .mi({\t/a/ID_op [4],open_n33672}),
    .sr(rst_pad),
    .f({_al_u1747_o,open_n33673}),
    .q({\t/a/EX_op [4],\t/a/ID_op [5]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0*D))"),
    //.LUTF1("0"),
    //.LUTG0("(C*B*A*~(1*D))"),
    //.LUTG1("A*~B*~C*D+A*B*~C*D+A*~B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000010000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0010101000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg6_b5|t/a/ex_mem/reg2_b5  (
    .a({_al_u2608_o,_al_u2608_o}),
    .b({_al_u1740_o,\t/a/risk_jump/n11_lutinv }),
    .c({\t/a/EX_op [5],\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({\t/a/risk_jump/n35_lutinv ,_al_u1740_o}),
    .e({\t/a/condition/n1_lutinv ,\t/a/EX_op [5]}),
    .mi({\t/a/ID_op [5],\t/a/EX_op [5]}),
    .sr(rst_pad),
    .f({_al_u2609_o,_al_u2615_o}),
    .q({\t/a/EX_op [5],\t/a/MEM_op [5]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUT1("(~(~C*~A)*~(D)*~(B)+~(~C*~A)*D*~(B)+~(~(~C*~A))*D*B+~(~C*~A)*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111100010),
    .INIT_LUT1(16'b1111111000110010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b11|t/a/id_ex/reg7_b30  (
    .a({_al_u2807_o,_al_u2807_o}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/memstraddress [11],\t/a/ID_memstraddr [30]}),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [11],\t/memstraddress [30]}),
    .mi({\t/a/ID_memstraddr [11],\t/a/ID_memstraddr [30]}),
    .sr(rst_pad),
    .f({_al_u2883_o,_al_u2829_o}),
    .q({\t/a/EX_memstraddr [11],\t/a/EX_memstraddr [30]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~C*~B*~D+A*~C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*~C*B*D+A*~C*B*D"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("A*~C*~B*~D+~A*C*~B*~D+A*C*~B*~D+A*~C*B*~D+~A*C*B*~D+A*C*B*~D+~A*~C*~B*D+A*~C*~B*D+~A*C*~B*D+A*C*~B*D+~A*~C*B*D+A*~C*B*D+~A*C*B*D+A*C*B*D"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100001010),
    .INIT_LUTF1(16'b1111000010101010),
    .INIT_LUTG0(16'b1111111111111010),
    .INIT_LUTG1(16'b1111000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b13|t/a/id_ex/reg7_b29  (
    .a({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/ID_memstraddr [13],\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/condition/n0_lutinv ,\t/memstraddress [29]}),
    .e({\t/memstraddress [13],\t/a/ID_memstraddr [29]}),
    .mi({\t/a/ID_memstraddr [13],\t/a/ID_memstraddr [29]}),
    .sr(rst_pad),
    .f({_al_u2878_o,_al_u2834_o}),
    .q({\t/a/EX_memstraddr [13],\t/a/EX_memstraddr [29]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("D*~A*~B*~C+D*~A*B*~C+~D*~A*~B*C+D*~A*~B*C+~D*~A*B*C+D*~A*B*C"),
    //.LUTF1("A*~D*~C*~B+A*D*~C*~B+A*~D*C*~B+A*D*C*~B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    //.LUTG0("D*~A*~B*~C+~D*A*~B*~C+D*A*~B*~C+D*~A*B*~C+~D*A*B*~C+D*A*B*~C+~D*~A*~B*C+D*~A*~B*C+~D*A*~B*C+D*A*~B*C+~D*~A*B*C+D*~A*B*C+~D*A*B*C+D*A*B*C"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010101010000),
    .INIT_LUTF1(16'b1110001011100010),
    .INIT_LUTG0(16'b1111111111111010),
    .INIT_LUTG1(16'b1111001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b14|t/a/id_ex/reg7_b26  (
    .a({_al_u2807_o,\t/a/condition/n0_lutinv }),
    .b({\t/a/condition/n0_lutinv ,open_n33725}),
    .c({\t/a/ID_memstraddr [14],\t/memstraddress [26]}),
    .clk(clock_pad),
    .d({open_n33727,_al_u2807_o}),
    .e({\t/memstraddress [14],\t/a/ID_memstraddr [26]}),
    .mi({\t/a/ID_memstraddr [14],\t/a/ID_memstraddr [26]}),
    .sr(rst_pad),
    .f({_al_u2875_o,_al_u2841_o}),
    .q({\t/a/EX_memstraddr [14],\t/a/EX_memstraddr [26]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUT1("(~(~C*~A)*~(D)*~(B)+~(~C*~A)*D*~(B)+~(~(~C*~A))*D*B+~(~C*~A)*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111100010),
    .INIT_LUT1(16'b1111111000110010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b15|t/a/id_ex/reg7_b25  (
    .a({_al_u2807_o,_al_u2807_o}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/memstraddress [15],\t/a/ID_memstraddr [25]}),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [15],\t/memstraddress [25]}),
    .mi({\t/a/ID_memstraddr [15],\t/a/ID_memstraddr [25]}),
    .sr(rst_pad),
    .f({_al_u2872_o,_al_u2844_o}),
    .q({\t/a/EX_memstraddr [15],\t/a/EX_memstraddr [25]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUT1("(~(~C*~A)*~(D)*~(B)+~(~C*~A)*D*~(B)+~(~(~C*~A))*D*B+~(~C*~A)*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111100010),
    .INIT_LUT1(16'b1111111000110010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b16|t/a/id_ex/reg7_b24  (
    .a({_al_u2807_o,_al_u2807_o}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/memstraddress [16],\t/a/ID_memstraddr [24]}),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [16],\t/memstraddress [24]}),
    .mi({\t/a/ID_memstraddr [16],\t/a/ID_memstraddr [24]}),
    .sr(rst_pad),
    .f({_al_u2869_o,_al_u2847_o}),
    .q({\t/a/EX_memstraddr [16],\t/a/EX_memstraddr [24]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("D*~B*~A*~C+D*~B*A*~C+~D*~B*~A*C+D*~B*~A*C+~D*~B*A*C+D*~B*A*C"),
    //.LUTF1("C*~B*~D*~A+~C*B*~D*~A+C*B*~D*~A+C*~B*D*~A+~C*B*D*~A+C*B*D*~A"),
    //.LUTG0("D*~B*~A*~C+~D*B*~A*~C+D*B*~A*~C+D*~B*A*~C+~D*B*A*~C+D*B*A*~C+~D*~B*~A*C+D*~B*~A*C+~D*B*~A*C+D*B*~A*C+~D*~B*A*C+D*~B*A*C+~D*B*A*C+D*B*A*C"),
    //.LUTG1("C*~B*~D*~A+~C*B*~D*~A+C*B*~D*~A+C*~B*D*~A+~C*B*D*~A+C*B*D*~A+~C*~B*~D*A+C*~B*~D*A+~C*B*~D*A+C*B*~D*A+~C*~B*D*A+C*~B*D*A+~C*B*D*A+C*B*D*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100110000),
    .INIT_LUTF1(16'b0101010001010100),
    .INIT_LUTG0(16'b1111111111111100),
    .INIT_LUTG1(16'b1111111011111110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b1|t/a/id_ex/reg7_b23  (
    .a({\t/a/condition/n0_lutinv ,open_n33771}),
    .b({\t/memstraddress [1],\t/a/condition/n0_lutinv }),
    .c({_al_u2807_o,\t/memstraddress [23]}),
    .clk(clock_pad),
    .d({open_n33773,_al_u2807_o}),
    .e({\t/a/ID_memstraddr [1],\t/a/ID_memstraddr [23]}),
    .mi({\t/a/ID_memstraddr [1],\t/a/ID_memstraddr [23]}),
    .sr(rst_pad),
    .f({_al_u2888_o,_al_u2850_o}),
    .q({\t/a/EX_memstraddr [1],\t/a/EX_memstraddr [23]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("A*~B*~D*~C+A*~B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*~B*D*C+A*~B*D*C"),
    //.LUTF1("C*~B*~D*~A+~C*B*~D*~A+C*B*~D*~A+C*~B*D*~A+~C*B*D*~A+C*B*D*~A"),
    //.LUTG0("A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    //.LUTG1("C*~B*~D*~A+~C*B*~D*~A+C*B*~D*~A+C*~B*D*~A+~C*B*D*~A+C*B*D*~A+~C*~B*~D*A+C*~B*~D*A+~C*B*~D*A+C*B*~D*A+~C*~B*D*A+C*~B*D*A+~C*B*D*A+C*B*D*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001000110010),
    .INIT_LUTF1(16'b0101010001010100),
    .INIT_LUTG0(16'b1111111011111110),
    .INIT_LUTG1(16'b1111111011111110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b2|t/a/id_ex/reg7_b20  (
    .a({\t/a/condition/n0_lutinv ,_al_u2807_o}),
    .b({\t/memstraddress [2],\t/a/condition/n0_lutinv }),
    .c({_al_u2807_o,\t/memstraddress [20]}),
    .clk(clock_pad),
    .e({\t/a/ID_memstraddr [2],\t/a/ID_memstraddr [20]}),
    .mi({\t/a/ID_memstraddr [2],\t/a/ID_memstraddr [20]}),
    .sr(rst_pad),
    .f({_al_u2860_o,_al_u2857_o}),
    .q({\t/a/EX_memstraddr [2],\t/a/EX_memstraddr [20]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1100110100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b0|t/a/id_ex/reg8_b9  (
    .a({_al_u994_o,_al_u333_o}),
    .b({_al_u333_o,_al_u343_o}),
    .c({_al_u1004_o,_al_u353_o}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [0],\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [0],\t/a/ID_read_dat1 [9]}),
    .q({\t/a/EX_regdat1 [0],\t/a/EX_regdat1 [9]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~D*~B)*~(C)*~(A)+(~D*~B)*C*~(A)+~((~D*~B))*C*A+(~D*~B)*C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1010000010110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b10|t/a/id_ex/reg8_b30  (
    .a({_al_u333_o,_al_u333_o}),
    .b({_al_u973_o,_al_u511_o}),
    .c({\t/a/reg_writedat [10],_al_u521_o}),
    .clk(clock_pad),
    .d({_al_u983_o,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [10],\t/a/ID_read_dat1 [30]}),
    .q({\t/a/EX_regdat1 [10],\t/a/EX_regdat1 [30]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~D*~A)*~(C)*~(B)+(~D*~A)*C*~(B)+~((~D*~A))*C*B+(~D*~A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1100000011010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b11|t/a/id_ex/reg8_b27  (
    .a({_al_u952_o,_al_u333_o}),
    .b({_al_u333_o,_al_u595_o}),
    .c({\t/a/reg_writedat [11],_al_u605_o}),
    .clk(clock_pad),
    .d({_al_u962_o,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [11],\t/a/ID_read_dat1 [27]}),
    .q({\t/a/EX_regdat1 [11],\t/a/EX_regdat1 [27]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~D*~A)*~(C)*~(B)+(~D*~A)*C*~(B)+~((~D*~A))*C*B+(~D*~A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1100000011010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b12|t/a/id_ex/reg8_b26  (
    .a({_al_u931_o,_al_u333_o}),
    .b({_al_u333_o,_al_u616_o}),
    .c({\t/a/reg_writedat [12],_al_u626_o}),
    .clk(clock_pad),
    .d({_al_u941_o,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [12],\t/a/ID_read_dat1 [26]}),
    .q({\t/a/EX_regdat1 [12],\t/a/EX_regdat1 [26]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~D*~B)*~(C)*~(A)+(~D*~B)*C*~(A)+~((~D*~B))*C*A+(~D*~B)*C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1010000010110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b13|t/a/id_ex/reg8_b23  (
    .a({_al_u333_o,_al_u333_o}),
    .b({_al_u910_o,_al_u679_o}),
    .c({\t/a/reg_writedat [13],_al_u689_o}),
    .clk(clock_pad),
    .d({_al_u920_o,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [13],\t/a/ID_read_dat1 [23]}),
    .q({\t/a/EX_regdat1 [13],\t/a/EX_regdat1 [23]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~C*~A)*~(D)*~(B)+(~C*~A)*D*~(B)+~((~C*~A))*D*B+(~C*~A)*D*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1100110100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b14|t/a/id_ex/reg8_b22  (
    .a({_al_u889_o,_al_u333_o}),
    .b({_al_u333_o,_al_u700_o}),
    .c({_al_u899_o,_al_u710_o}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [14],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [14],\t/a/ID_read_dat1 [22]}),
    .q({\t/a/EX_regdat1 [14],\t/a/EX_regdat1 [22]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~D*~B)*~(C)*~(A)+(~D*~B)*C*~(A)+~((~D*~B))*C*A+(~D*~B)*C*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1010000010110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b15|t/a/id_ex/reg8_b19  (
    .a({_al_u333_o,_al_u333_o}),
    .b({_al_u868_o,_al_u784_o}),
    .c({\t/a/reg_writedat [15],_al_u794_o}),
    .clk(clock_pad),
    .d({_al_u878_o,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [15],\t/a/ID_read_dat1 [19]}),
    .q({\t/a/EX_regdat1 [15],\t/a/EX_regdat1 [19]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("~A*B*~D*~C+~A*B*D*~C+~A*B*~D*C+~A*B*D*C"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("~A*~B*D*~C+~A*B*D*~C+~A*~B*D*C+~A*B*D*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0100010001000100),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0101010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b0|t/a/id_ex/reg2_b0  (
    .a({\t/a/if_id/n9 ,\t/a/condition/n5 [5]}),
    .b({\t/busarbitration/instruction [25],\t/a/condition/n0_lutinv }),
    .c({open_n33919,\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({i_data[25],\t/a/condition/sel1/B2 }),
    .e({\t/busarbitration/n3 ,\t/a/ID_fun7 [0]}),
    .mi({open_n33922,\t/a/ID_fun7 [0]}),
    .sr(rst_pad),
    .f({open_n33934,\t/a/ID_jump_addr [5]}),
    .q({\t/a/ID_fun7 [0],\t/a/EX_fun7 [0]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("~C*A*~B*~D+C*A*~B*~D+~C*A*B*~D+C*A*B*~D+~C*~A*B*D+C*~A*B*D+~C*A*B*D+C*A*B*D"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b1100110010101010),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b1|t/a/id_ex/reg2_b1  (
    .a({\t/busarbitration/instruction [26],\t/a/condition/n5 [6]}),
    .b({i_data[26],\t/a/condition/n0_lutinv }),
    .c({open_n33938,\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,\t/a/condition/sel1/B2 }),
    .e({\t/a/if_id/n9 ,\t/a/ID_fun7 [1]}),
    .mi({open_n33941,\t/a/ID_fun7 [1]}),
    .sr(rst_pad),
    .f({open_n33953,\t/a/ID_jump_addr [6]}),
    .q({\t/a/ID_fun7 [1],\t/a/EX_fun7 [1]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b1110001011100010),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b2|t/a/id_ex/reg2_b2  (
    .a({\t/busarbitration/instruction [27],\t/a/condition/n5 [7]}),
    .b({\t/busarbitration/n3 ,\t/a/condition/n0_lutinv }),
    .c({i_data[27],\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({open_n33958,\t/a/condition/sel1/B2 }),
    .e({\t/a/if_id/n9 ,\t/a/ID_fun7 [2]}),
    .mi({open_n33960,\t/a/ID_fun7 [2]}),
    .sr(rst_pad),
    .f({open_n33972,\t/a/ID_jump_addr [7]}),
    .q({\t/a/ID_fun7 [2],\t/a/EX_fun7 [2]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("~D*~A*C*~B+D*~A*C*~B+~D*A*~C*B+D*A*~C*B+~D*~A*C*B+D*~A*C*B+~D*A*C*B+D*A*C*B"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b1101100011011000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b3|t/a/id_ex/reg2_b3  (
    .a({\t/busarbitration/n3 ,\t/a/condition/n5 [8]}),
    .b({i_data[28],\t/a/condition/n0_lutinv }),
    .c({\t/busarbitration/instruction [28],\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({open_n33977,\t/a/condition/sel1/B2 }),
    .e({\t/a/if_id/n9 ,\t/a/ID_fun7 [3]}),
    .mi({open_n33979,\t/a/ID_fun7 [3]}),
    .sr(rst_pad),
    .f({open_n33991,\t/a/ID_jump_addr [8]}),
    .q({\t/a/ID_fun7 [3],\t/a/EX_fun7 [3]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("C*~A*~B*~D+C*A*~B*~D+C*~A*B*~D+C*A*B*~D+~C*A*~B*D+C*A*~B*D+~C*A*B*D+C*A*B*D"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b1010101011110000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b4|t/a/id_ex/reg2_b4  (
    .a({i_data[29],\t/a/condition/n5 [9]}),
    .b({open_n33995,\t/a/condition/n0_lutinv }),
    .c({\t/busarbitration/instruction [29],\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,\t/a/condition/sel1/B2 }),
    .e({\t/a/if_id/n9 ,\t/a/ID_fun7 [4]}),
    .mi({open_n33998,\t/a/ID_fun7 [4]}),
    .sr(rst_pad),
    .f({open_n34010,\t/a/ID_jump_addr [9]}),
    .q({\t/a/ID_fun7 [4],\t/a/EX_fun7 [4]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b1100110010101010),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b5|t/a/id_ex/reg2_b5  (
    .a({\t/busarbitration/instruction [30],\t/a/condition/n5 [10]}),
    .b({i_data[30],\t/a/condition/n0_lutinv }),
    .c({open_n34014,\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,\t/a/condition/sel1/B2 }),
    .e({\t/a/if_id/n9 ,\t/a/ID_fun7 [5]}),
    .mi({open_n34017,\t/a/ID_fun7 [5]}),
    .sr(rst_pad),
    .f({open_n34029,\t/a/ID_jump_addr [10]}),
    .q({\t/a/ID_fun7 [5],\t/a/EX_fun7 [5]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)"),
    //.LUTF1("B*~A*~C*~D+B*A*~C*~D+B*~A*~C*D+B*A*~C*D"),
    //.LUTG0("(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)"),
    //.LUTG1("B*~A*~C*~D+B*A*~C*~D+~B*~A*C*~D+B*~A*C*~D+~B*A*C*~D+B*A*C*~D+B*~A*~C*D+B*A*~C*D+~B*~A*C*D+B*~A*C*D+~B*A*C*D+B*A*C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010110100000),
    .INIT_LUTF1(16'b0000110000001100),
    .INIT_LUTG0(16'b1111010110100000),
    .INIT_LUTG1(16'b1111110011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b10|t/a/if_id/reg5_b8  (
    .a({open_n34033,\t/busarbitration/n3_placeOpt_5 }),
    .b({\t/a/MEM_aludat [10],open_n34034}),
    .c({\t/busarbitration/n3_placeOpt_5 ,\t/memstraddress [8]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({open_n34035,\t/a/MEM_aludat [8]}),
    .e({\t/memstraddress [10],open_n34036}),
    .mi({\t/memstraddress [10],\t/memstraddress [8]}),
    .sr(rst_pad),
    .f({addr[10],addr[8]}),
    .q({\t/a/ID_memstraddr [10],\t/a/ID_memstraddr [8]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)"),
    //.LUTF1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTG0("(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101011110000),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b1010101011110000),
    .INIT_LUTG1(16'b1111111111001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b11|t/a/if_id/reg5_b30  (
    .a({open_n34052,\t/memstraddress [30]}),
    .b({\t/a/MEM_aludat [11],open_n34053}),
    .c({open_n34054,\t/a/MEM_aludat [30]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/busarbitration/n3_placeOpt_1 ,\t/busarbitration/n3_placeOpt_1 }),
    .e({\t/memstraddress [11],open_n34055}),
    .mi({\t/memstraddress [11],\t/memstraddress [30]}),
    .sr(rst_pad),
    .f({addr[11],addr[30]}),
    .q({\t/a/ID_memstraddr [11],\t/a/ID_memstraddr [30]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)"),
    //.LUT1("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101011001100),
    .INIT_LUT1(16'b1101100011011000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b12|t/a/if_id/reg5_b28  (
    .a({\t/busarbitration/n3_placeOpt_1 ,\t/memstraddress [28]}),
    .b({\t/memstraddress [12],\t/a/MEM_aludat [28]}),
    .c({\t/a/MEM_aludat [12],open_n34071}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({open_n34072,\t/busarbitration/n3_placeOpt_1 }),
    .mi({\t/memstraddress [12],\t/memstraddress [28]}),
    .sr(rst_pad),
    .f({addr[12],addr[28]}),
    .q({\t/a/ID_memstraddr [12],\t/a/ID_memstraddr [28]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("B*~A*~D*~C+B*A*~D*~C+B*~A*~D*C+B*A*~D*C"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("B*~A*~D*~C+B*A*~D*~C+~B*~A*D*~C+B*~A*D*~C+~B*A*D*~C+B*A*D*~C+B*~A*~D*C+B*A*~D*C+~B*~A*D*C+B*~A*D*C+~B*A*D*C+B*A*D*C"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111111111001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b13|t/a/if_id/reg5_b27  (
    .b({\t/a/MEM_aludat [13],\t/a/MEM_aludat [27]}),
    .c({open_n34088,\t/memstraddress [27]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/busarbitration/n3_placeOpt_1 ,\t/busarbitration/n3_placeOpt_1 }),
    .e({\t/memstraddress [13],open_n34089}),
    .mi({\t/memstraddress [13],\t/memstraddress [27]}),
    .sr(rst_pad),
    .f({addr[13],addr[27]}),
    .q({\t/a/ID_memstraddr [13],\t/a/ID_memstraddr [27]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A)"),
    //.LUT1("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010110100000),
    .INIT_LUT1(16'b1011100010111000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b14|t/a/if_id/reg5_b25  (
    .a({\t/memstraddress [14],\t/busarbitration/n3_placeOpt_1 }),
    .b({\t/busarbitration/n3_placeOpt_1 ,open_n34105}),
    .c({\t/a/MEM_aludat [14],\t/memstraddress [25]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({open_n34106,\t/a/MEM_aludat [25]}),
    .mi({\t/memstraddress [14],\t/memstraddress [25]}),
    .sr(rst_pad),
    .f({addr[14],addr[25]}),
    .q({\t/a/ID_memstraddr [14],\t/a/ID_memstraddr [25]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    //.LUTF1("~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011001100),
    .INIT_LUTF1(16'b1111111100000000),
    .INIT_LUTG0(16'b1111111111001100),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b15|t/a/if_id/reg5_b23  (
    .a({\t/memstraddress [15],open_n34120}),
    .b({open_n34121,\t/a/MEM_aludat [23]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [15],\t/busarbitration/n3_placeOpt_1 }),
    .e({\t/busarbitration/n3_placeOpt_1 ,\t/memstraddress [23]}),
    .mi({\t/memstraddress [15],\t/memstraddress [23]}),
    .sr(rst_pad),
    .f({addr[15],addr[23]}),
    .q({\t/a/ID_memstraddr [15],\t/a/ID_memstraddr [23]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    //.LUT1("(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010110010101100),
    .INIT_LUT1(16'b1111001111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b16|t/a/if_id/reg5_b21  (
    .a({open_n34139,\t/memstraddress [21]}),
    .b({\t/busarbitration/n3_placeOpt_1 ,\t/a/MEM_aludat [21]}),
    .c({\t/memstraddress [16],\t/busarbitration/n3_placeOpt_1 }),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [16],open_n34140}),
    .mi({\t/memstraddress [16],\t/memstraddress [21]}),
    .sr(rst_pad),
    .f({addr[16],addr[21]}),
    .q({\t/a/ID_memstraddr [16],\t/a/ID_memstraddr [21]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    //.LUT1("(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010110010101100),
    .INIT_LUT1(16'b1111110000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b17|t/a/if_id/reg5_b20  (
    .a({open_n34154,\t/memstraddress [20]}),
    .b({\t/busarbitration/n3 ,\t/a/MEM_aludat [20]}),
    .c({\t/a/MEM_aludat [17],\t/busarbitration/n3 }),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/memstraddress [17],open_n34155}),
    .mi({\t/memstraddress [17],\t/memstraddress [20]}),
    .sr(rst_pad),
    .f({addr[17],addr[20]}),
    .q({\t/a/ID_memstraddr [17],\t/a/ID_memstraddr [20]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u11_al_u2955  (
    .a({\t/memstraddress [13],\t/memstraddress [11]}),
    .b({\t/memstraddress [14],\t/memstraddress [12]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [13],\t/a/IF_skip_addr [11]}),
    .e({\t/a/IF_skip_addr [14],\t/a/IF_skip_addr [12]}),
    .fci(\t/a/instr/add0/c11 ),
    .f({\t/a/instr/n12 [13],\t/a/instr/n12 [11]}),
    .fco(\t/a/instr/add0/c15 ),
    .fx({\t/a/instr/n12 [14],\t/a/instr/n12 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u15_al_u2956  (
    .a({\t/memstraddress [17],\t/memstraddress [15]}),
    .b({\t/memstraddress [18],\t/memstraddress [16]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [17],\t/a/IF_skip_addr [15]}),
    .e({\t/a/IF_skip_addr [18],\t/a/IF_skip_addr [16]}),
    .fci(\t/a/instr/add0/c15 ),
    .f({\t/a/instr/n12 [17],\t/a/instr/n12 [15]}),
    .fco(\t/a/instr/add0/c19 ),
    .fx({\t/a/instr/n12 [18],\t/a/instr/n12 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u19_al_u2957  (
    .a({\t/memstraddress [21],\t/memstraddress [19]}),
    .b({\t/memstraddress [22],\t/memstraddress [20]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [21],\t/a/IF_skip_addr [19]}),
    .e({\t/a/IF_skip_addr [22],\t/a/IF_skip_addr [20]}),
    .fci(\t/a/instr/add0/c19 ),
    .f({\t/a/instr/n12 [21],\t/a/instr/n12 [19]}),
    .fco(\t/a/instr/add0/c23 ),
    .fx({\t/a/instr/n12 [22],\t/a/instr/n12 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u23_al_u2958  (
    .a({\t/memstraddress [25],\t/memstraddress [23]}),
    .b({\t/memstraddress [26],\t/memstraddress [24]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [25],\t/a/IF_skip_addr [23]}),
    .e({\t/a/IF_skip_addr [26],\t/a/IF_skip_addr [24]}),
    .fci(\t/a/instr/add0/c23 ),
    .f({\t/a/instr/n12 [25],\t/a/instr/n12 [23]}),
    .fco(\t/a/instr/add0/c27 ),
    .fx({\t/a/instr/n12 [26],\t/a/instr/n12 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u27_al_u2959  (
    .a({\t/memstraddress [29],\t/memstraddress [27]}),
    .b({\t/memstraddress [30],\t/memstraddress [28]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [29],\t/a/IF_skip_addr [27]}),
    .e({\t/a/IF_skip_addr [30],\t/a/IF_skip_addr [28]}),
    .fci(\t/a/instr/add0/c27 ),
    .f({\t/a/instr/n12 [29],\t/a/instr/n12 [27]}),
    .fco(\t/a/instr/add0/c31 ),
    .fx({\t/a/instr/n12 [30],\t/a/instr/n12 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u31_al_u2960  (
    .a({open_n34259,\t/memstraddress [31]}),
    .c(2'b00),
    .d({open_n34264,\t/a/IF_skip_addr [31]}),
    .fci(\t/a/instr/add0/c31 ),
    .f({open_n34281,\t/a/instr/n12 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u3_al_u2953  (
    .a({\t/memstraddress [5],\t/memstraddress [3]}),
    .b({\t/memstraddress [6],\t/memstraddress [4]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [5],\t/a/IF_skip_addr [3]}),
    .e({\t/a/IF_skip_addr [6],\t/a/IF_skip_addr [4]}),
    .fci(\t/a/instr/add0/c3 ),
    .f({\t/a/instr/n12 [5],\t/a/instr/n12 [3]}),
    .fco(\t/a/instr/add0/c7 ),
    .fx({\t/a/instr/n12 [6],\t/a/instr/n12 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u7_al_u2954  (
    .a({\t/memstraddress [9],\t/memstraddress [7]}),
    .b({\t/memstraddress [10],\t/memstraddress [8]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [9],\t/a/IF_skip_addr [7]}),
    .e({\t/a/IF_skip_addr [10],\t/a/IF_skip_addr [8]}),
    .fci(\t/a/instr/add0/c7 ),
    .f({\t/a/instr/n12 [9],\t/a/instr/n12 [7]}),
    .fco(\t/a/instr/add0/c11 ),
    .fx({\t/a/instr/n12 [10],\t/a/instr/n12 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/add0/ucin_al_u2952  (
    .a({\t/memstraddress [1],1'b0}),
    .b({\t/memstraddress [2],\t/memstraddress [0]}),
    .c(2'b00),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/a/IF_skip_addr [1],1'b1}),
    .e({\t/a/IF_skip_addr [2],1'b0}),
    .mi({open_n34324,\t/memstraddress [0]}),
    .sr(rst_pad),
    .f({\t/a/instr/n12 [1],open_n34336}),
    .fco(\t/a/instr/add0/c3 ),
    .fx({\t/a/instr/n12 [2],\t/a/instr/n12 [0]}),
    .q({open_n34337,\t/a/ID_memstraddr [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u11_al_u2972  (
    .a({\t/memstraddress [15],\t/memstraddress [13]}),
    .b({\t/memstraddress [16],\t/memstraddress [14]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c11 ),
    .f({\t/a/instr/n16 [13],\t/a/instr/n16 [11]}),
    .fco(\t/a/instr/add2/c15 ),
    .fx({\t/a/instr/n16 [14],\t/a/instr/n16 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u15_al_u2973  (
    .a({\t/memstraddress [19],\t/memstraddress [17]}),
    .b({\t/memstraddress [20],\t/memstraddress [18]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c15 ),
    .f({\t/a/instr/n16 [17],\t/a/instr/n16 [15]}),
    .fco(\t/a/instr/add2/c19 ),
    .fx({\t/a/instr/n16 [18],\t/a/instr/n16 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u19_al_u2974  (
    .a({\t/memstraddress [23],\t/memstraddress [21]}),
    .b({\t/memstraddress [24],\t/memstraddress [22]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c19 ),
    .f({\t/a/instr/n16 [21],\t/a/instr/n16 [19]}),
    .fco(\t/a/instr/add2/c23 ),
    .fx({\t/a/instr/n16 [22],\t/a/instr/n16 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u23_al_u2975  (
    .a({\t/memstraddress [27],\t/memstraddress [25]}),
    .b({\t/memstraddress [28],\t/memstraddress [26]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c23 ),
    .f({\t/a/instr/n16 [25],\t/a/instr/n16 [23]}),
    .fco(\t/a/instr/add2/c27 ),
    .fx({\t/a/instr/n16 [26],\t/a/instr/n16 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u27_al_u2976  (
    .a({\t/memstraddress [31],\t/memstraddress [29]}),
    .b({open_n34410,\t/memstraddress [30]}),
    .c(2'b00),
    .d(2'b00),
    .e({open_n34413,1'b0}),
    .fci(\t/a/instr/add2/c27 ),
    .f({\t/a/instr/n16 [29],\t/a/instr/n16 [27]}),
    .fx({open_n34429,\t/a/instr/n16 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u3_al_u2970  (
    .a({\t/memstraddress [7],\t/memstraddress [5]}),
    .b({\t/memstraddress [8],\t/memstraddress [6]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c3 ),
    .f({\t/a/instr/n16 [5],\t/a/instr/n16 [3]}),
    .fco(\t/a/instr/add2/c7 ),
    .fx({\t/a/instr/n16 [6],\t/a/instr/n16 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u7_al_u2971  (
    .a({\t/memstraddress [11],\t/memstraddress [9]}),
    .b({\t/memstraddress [12],\t/memstraddress [10]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c7 ),
    .f({\t/a/instr/n16 [9],\t/a/instr/n16 [7]}),
    .fco(\t/a/instr/add2/c11 ),
    .fx({\t/a/instr/n16 [10],\t/a/instr/n16 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/add2/ucin_al_u2969  (
    .a({\t/memstraddress [3],1'b0}),
    .b({\t/memstraddress [4],\t/memstraddress [2]}),
    .c(2'b00),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d(2'b01),
    .e(2'b01),
    .mi(\t/memstraddress [4:3]),
    .sr(rst_pad),
    .f({\t/a/instr/n16 [1],open_n34480}),
    .fco(\t/a/instr/add2/c3 ),
    .fx({\t/a/instr/n16 [2],\t/a/instr/n16 [0]}),
    .q(\t/a/ID_memstraddr [4:3]));
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b0  (
    .a({_al_u2890_o,_al_u2890_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [0],\t/a/ID_memstraddr [0]}),
    .mi({open_n34492,\t/memstraddress [0]}),
    .sr(rst_pad),
    .q({open_n34498,\t/memstraddress [0]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b1  (
    .a({_al_u2887_o,_al_u2887_o}),
    .b({\t/a/instr/n12 [1],\t/a/instr/n12 [1]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2888_o,_al_u2888_o}),
    .mi({open_n34510,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34516,\t/memstraddress [1]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b10  (
    .a({_al_u2885_o,_al_u2885_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [10],\t/a/ID_memstraddr [10]}),
    .mi({open_n34528,\t/memstraddress [10]}),
    .sr(rst_pad),
    .q({open_n34534,\t/memstraddress [10]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b11  (
    .a({_al_u2882_o,_al_u2882_o}),
    .b({\t/a/instr/n12 [11],\t/a/instr/n12 [11]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2883_o,_al_u2883_o}),
    .mi({open_n34546,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34552,\t/memstraddress [11]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b12  (
    .a({_al_u2880_o,_al_u2880_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [12],\t/a/ID_memstraddr [12]}),
    .mi({open_n34564,\t/memstraddress [12]}),
    .sr(rst_pad),
    .q({open_n34570,\t/memstraddress [12]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b13  (
    .a({_al_u2877_o,_al_u2877_o}),
    .b({\t/a/instr/n12 [13],\t/a/instr/n12 [13]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2878_o,_al_u2878_o}),
    .mi({open_n34582,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34588,\t/memstraddress [13]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b14  (
    .a({_al_u2874_o,_al_u2874_o}),
    .b({\t/a/instr/n12 [14],\t/a/instr/n12 [14]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2875_o,_al_u2875_o}),
    .mi({open_n34600,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34606,\t/memstraddress [14]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b15  (
    .a({_al_u2871_o,_al_u2871_o}),
    .b({\t/a/instr/n12 [15],\t/a/instr/n12 [15]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2872_o,_al_u2872_o}),
    .mi({open_n34618,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34624,\t/memstraddress [15]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b16  (
    .a({_al_u2868_o,_al_u2868_o}),
    .b({\t/a/instr/n12 [16],\t/a/instr/n12 [16]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2869_o,_al_u2869_o}),
    .mi({open_n34636,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34642,\t/memstraddress [16]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b17  (
    .a({_al_u2866_o,_al_u2866_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [17],\t/a/ID_memstraddr [17]}),
    .mi({open_n34654,\t/memstraddress [17]}),
    .sr(rst_pad),
    .q({open_n34660,\t/memstraddress [17]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b18  (
    .a({_al_u2864_o,_al_u2864_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [18],\t/a/ID_memstraddr [18]}),
    .mi({open_n34672,\t/memstraddress [18]}),
    .sr(rst_pad),
    .q({open_n34678,\t/memstraddress [18]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b19  (
    .a({_al_u2862_o,_al_u2862_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [19],\t/a/ID_memstraddr [19]}),
    .mi({open_n34690,\t/memstraddress [19]}),
    .sr(rst_pad),
    .q({open_n34696,\t/memstraddress [19]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("SET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b2  (
    .a({_al_u2859_o,_al_u2859_o}),
    .b({\t/a/instr/n12 [2],\t/a/instr/n12 [2]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2860_o,_al_u2860_o}),
    .mi({open_n34708,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34714,\t/memstraddress [2]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b20  (
    .a({_al_u2856_o,_al_u2856_o}),
    .b({\t/a/instr/n12 [20],\t/a/instr/n12 [20]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2857_o,_al_u2857_o}),
    .mi({open_n34726,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34732,\t/memstraddress [20]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b21  (
    .a({_al_u2854_o,_al_u2854_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [21],\t/a/ID_memstraddr [21]}),
    .mi({open_n34744,\t/memstraddress [21]}),
    .sr(rst_pad),
    .q({open_n34750,\t/memstraddress [21]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b22  (
    .a({_al_u2852_o,_al_u2852_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [22],\t/a/ID_memstraddr [22]}),
    .mi({open_n34762,\t/memstraddress [22]}),
    .sr(rst_pad),
    .q({open_n34768,\t/memstraddress [22]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b23  (
    .a({_al_u2849_o,_al_u2849_o}),
    .b({\t/a/instr/n12 [23],\t/a/instr/n12 [23]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2850_o,_al_u2850_o}),
    .mi({open_n34780,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34786,\t/memstraddress [23]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b24  (
    .a({_al_u2846_o,_al_u2846_o}),
    .b({\t/a/instr/n12 [24],\t/a/instr/n12 [24]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2847_o,_al_u2847_o}),
    .mi({open_n34798,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34804,\t/memstraddress [24]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b25  (
    .a({_al_u2843_o,_al_u2843_o}),
    .b({\t/a/instr/n12 [25],\t/a/instr/n12 [25]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2844_o,_al_u2844_o}),
    .mi({open_n34816,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34822,\t/memstraddress [25]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b26  (
    .a({_al_u2840_o,_al_u2840_o}),
    .b({\t/a/instr/n12 [26],\t/a/instr/n12 [26]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2841_o,_al_u2841_o}),
    .mi({open_n34834,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34840,\t/memstraddress [26]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b27  (
    .a({_al_u2838_o,_al_u2838_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [27],\t/a/ID_memstraddr [27]}),
    .mi({open_n34852,\t/memstraddress [27]}),
    .sr(rst_pad),
    .q({open_n34858,\t/memstraddress [27]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b28  (
    .a({_al_u2836_o,_al_u2836_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [28],\t/a/ID_memstraddr [28]}),
    .mi({open_n34870,\t/memstraddress [28]}),
    .sr(rst_pad),
    .q({open_n34876,\t/memstraddress [28]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b29  (
    .a({_al_u2833_o,_al_u2833_o}),
    .b({\t/a/instr/n12 [29],\t/a/instr/n12 [29]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2834_o,_al_u2834_o}),
    .mi({open_n34888,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34894,\t/memstraddress [29]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b3  (
    .a({_al_u2831_o,_al_u2831_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [3],\t/a/ID_memstraddr [3]}),
    .mi({open_n34906,\t/memstraddress [3]}),
    .sr(rst_pad),
    .q({open_n34912,\t/memstraddress [3]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b30  (
    .a({_al_u2828_o,_al_u2828_o}),
    .b({\t/a/instr/n12 [30],\t/a/instr/n12 [30]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2829_o,_al_u2829_o}),
    .mi({open_n34924,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34930,\t/memstraddress [30]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b31  (
    .a({_al_u2826_o,_al_u2826_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [31],\t/a/ID_memstraddr [31]}),
    .mi({open_n34942,\t/memstraddress [31]}),
    .sr(rst_pad),
    .q({open_n34948,\t/memstraddress [31]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b4  (
    .a({_al_u2824_o,_al_u2824_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [4],\t/a/ID_memstraddr [4]}),
    .mi({open_n34960,\t/memstraddress [4]}),
    .sr(rst_pad),
    .q({open_n34966,\t/memstraddress [4]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b5  (
    .a({_al_u2821_o,_al_u2821_o}),
    .b({\t/a/instr/n12 [5],\t/a/instr/n12 [5]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2822_o,_al_u2822_o}),
    .mi({open_n34978,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n34984,\t/memstraddress [5]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b6  (
    .a({_al_u2819_o,_al_u2819_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [6],\t/a/ID_memstraddr [6]}),
    .mi({open_n34996,\t/memstraddress [6]}),
    .sr(rst_pad),
    .q({open_n35002,\t/memstraddress [6]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b7  (
    .a({_al_u2817_o,_al_u2817_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [7],\t/a/ID_memstraddr [7]}),
    .mi({open_n35014,\t/memstraddress [7]}),
    .sr(rst_pad),
    .q({open_n35020,\t/memstraddress [7]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b8  (
    .a({_al_u2814_o,_al_u2814_o}),
    .b({\t/a/instr/n12 [8],\t/a/instr/n12 [8]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2815_o,_al_u2815_o}),
    .mi({open_n35032,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n35038,\t/memstraddress [8]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b9  (
    .a({_al_u2811_o,_al_u2811_o}),
    .b({\t/a/instr/n12 [9],\t/a/instr/n12 [9]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2812_o,_al_u2812_o}),
    .mi({open_n35050,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n35056,\t/memstraddress [9]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~((0*~C))*~(B)+D*(0*~C)*~(B)+~(D)*(0*~C)*B+D*(0*~C)*B))"),
    //.LUT1("~(~B*~(D*~((1*~C))*~(A)+D*(1*~C)*~(A)+~(D)*(1*~C)*A+D*(1*~C)*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1101111111001110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b10  (
    .a({\t/busarbitration/mux5_b0_sel_is_3_o ,_al_u1902_o}),
    .b({_al_u1902_o,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .c({_al_u1903_o,_al_u1903_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [10],\t/a/MEM_aludat [10]}),
    .mi({open_n35068,i_data[10]}),
    .sr(rst_pad),
    .q({open_n35074,\t/a/reg_writedat [10]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*~C))"),
    //.LUT1("~(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111111101110),
    .INIT_LUT1(16'b1111111011011100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b11|t/a/mem_wb/reg0_b9  (
    .a({\t/busarbitration/mux5_b0_sel_is_3_o ,_al_u1902_o}),
    .b({_al_u1902_o,_al_u1904_o}),
    .c({\t/a/MEM_aludat [11],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({_al_u1940_o,\t/a/MEM_aludat [9]}),
    .sr(rst_pad),
    .q({\t/a/reg_writedat [11],\t/a/reg_writedat [9]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~((0*~C))*~(B)+D*(0*~C)*~(B)+~(D)*(0*~C)*B+D*(0*~C)*B))"),
    //.LUT1("~(~A*~(D*~((1*~C))*~(B)+D*(1*~C)*~(B)+~(D)*(1*~C)*B+D*(1*~C)*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1011111110101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b12  (
    .a({_al_u1902_o,_al_u1902_o}),
    .b({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .c({_al_u1903_o,_al_u1903_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [12],\t/a/MEM_aludat [12]}),
    .mi({open_n35104,i_data[12]}),
    .sr(rst_pad),
    .q({open_n35110,\t/a/reg_writedat [12]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~((0*~C))*~(B)+D*(0*~C)*~(B)+~(D)*(0*~C)*B+D*(0*~C)*B))"),
    //.LUT1("~(~B*~(D*~((1*~C))*~(A)+D*(1*~C)*~(A)+~(D)*(1*~C)*A+D*(1*~C)*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1101111111001110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b13  (
    .a({\t/busarbitration/mux5_b0_sel_is_3_o ,_al_u1902_o}),
    .b({_al_u1902_o,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .c({_al_u1903_o,_al_u1903_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [13],\t/a/MEM_aludat [13]}),
    .mi({open_n35122,i_data[13]}),
    .sr(rst_pad),
    .q({open_n35128,\t/a/reg_writedat [13]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~((0*~C))*~(B)+D*(0*~C)*~(B)+~(D)*(0*~C)*B+D*(0*~C)*B))"),
    //.LUT1("~(~B*~(C*~((1*~D))*~(A)+C*(1*~D)*~(A)+~(C)*(1*~D)*A+C*(1*~D)*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1101110011111110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b14  (
    .a({\t/busarbitration/mux5_b0_sel_is_3_o ,_al_u1902_o}),
    .b({_al_u1902_o,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .c({\t/a/MEM_aludat [14],_al_u1903_o}),
    .clk(clock_pad),
    .d({_al_u1903_o,\t/a/MEM_aludat [14]}),
    .mi({open_n35140,i_data[14]}),
    .sr(rst_pad),
    .q({open_n35146,\t/a/reg_writedat [14]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(B*~C)*~(1*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1111111110101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b16  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({\t/a/MEM_aludat [16],_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({_al_u1918_o,\t/a/MEM_aludat [16]}),
    .mi({open_n35158,i_data[16]}),
    .sr(rst_pad),
    .q({open_n35164,\t/a/reg_writedat [16]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~B*~(D*~C)*~(1*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b17  (
    .a({_al_u1918_o,_al_u1917_o}),
    .b({_al_u1917_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [17],\t/a/MEM_aludat [17]}),
    .mi({open_n35176,i_data[17]}),
    .sr(rst_pad),
    .q({open_n35182,\t/a/reg_writedat [17]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~B*~(C*~D)*~(1*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111011111110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b18  (
    .a({_al_u1918_o,_al_u1917_o}),
    .b({_al_u1917_o,_al_u1918_o}),
    .c({\t/a/MEM_aludat [18],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/a/MEM_aludat [18]}),
    .mi({open_n35194,i_data[18]}),
    .sr(rst_pad),
    .q({open_n35200,\t/a/reg_writedat [18]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~B*~(D*~C)*~(1*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b19  (
    .a({_al_u1918_o,_al_u1917_o}),
    .b({_al_u1917_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [19],\t/a/MEM_aludat [19]}),
    .mi({open_n35212,i_data[19]}),
    .sr(rst_pad),
    .q({open_n35218,\t/a/reg_writedat [19]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~B*~(A*~D)*~(1*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1111110011111110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b20  (
    .a({\t/a/MEM_aludat [20],_al_u1917_o}),
    .b({_al_u1917_o,_al_u1918_o}),
    .c({_al_u1918_o,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/a/MEM_aludat [20]}),
    .mi({open_n35230,i_data[20]}),
    .sr(rst_pad),
    .q({open_n35236,\t/a/reg_writedat [20]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b21  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [21],\t/a/MEM_aludat [21]}),
    .mi({open_n35248,i_data[21]}),
    .sr(rst_pad),
    .q({open_n35254,\t/a/reg_writedat [21]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~B*~(D*~C)*~(1*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b22  (
    .a({_al_u1918_o,_al_u1917_o}),
    .b({_al_u1917_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [22],\t/a/MEM_aludat [22]}),
    .mi({open_n35266,i_data[22]}),
    .sr(rst_pad),
    .q({open_n35272,\t/a/reg_writedat [22]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(B*~C)*~(1*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1111111110101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b23  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({\t/a/MEM_aludat [23],_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({_al_u1918_o,\t/a/MEM_aludat [23]}),
    .mi({open_n35284,i_data[23]}),
    .sr(rst_pad),
    .q({open_n35290,\t/a/reg_writedat [23]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~B*~(A*~C)*~(1*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1111111111001110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b24  (
    .a({\t/a/MEM_aludat [24],_al_u1917_o}),
    .b({_al_u1917_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({_al_u1918_o,\t/a/MEM_aludat [24]}),
    .mi({open_n35302,i_data[24]}),
    .sr(rst_pad),
    .q({open_n35308,\t/a/reg_writedat [24]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(B*~C)*~(1*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1111111110101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b25  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({\t/a/MEM_aludat [25],_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({_al_u1918_o,\t/a/MEM_aludat [25]}),
    .mi({open_n35320,i_data[25]}),
    .sr(rst_pad),
    .q({open_n35326,\t/a/reg_writedat [25]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~B*~(C*~D)*~(1*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111011111110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b26  (
    .a({_al_u1918_o,_al_u1917_o}),
    .b({_al_u1917_o,_al_u1918_o}),
    .c({\t/a/MEM_aludat [26],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/a/MEM_aludat [26]}),
    .mi({open_n35338,i_data[26]}),
    .sr(rst_pad),
    .q({open_n35344,\t/a/reg_writedat [26]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~B*~(D*~C)*~(1*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b27  (
    .a({_al_u1918_o,_al_u1917_o}),
    .b({_al_u1917_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [27],\t/a/MEM_aludat [27]}),
    .mi({open_n35356,i_data[27]}),
    .sr(rst_pad),
    .q({open_n35362,\t/a/reg_writedat [27]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(B*~C)*~(1*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1111111110101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b28  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({\t/a/MEM_aludat [28],_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({_al_u1918_o,\t/a/MEM_aludat [28]}),
    .mi({open_n35374,i_data[28]}),
    .sr(rst_pad),
    .q({open_n35380,\t/a/reg_writedat [28]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~B*~(D*~C)*~(1*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b29  (
    .a({_al_u1918_o,_al_u1917_o}),
    .b({_al_u1917_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [29],\t/a/MEM_aludat [29]}),
    .mi({open_n35392,i_data[29]}),
    .sr(rst_pad),
    .q({open_n35398,\t/a/reg_writedat [29]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~B*~(D*~C)*~(1*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b30  (
    .a({_al_u1918_o,_al_u1917_o}),
    .b({_al_u1917_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [30],\t/a/MEM_aludat [30]}),
    .mi({open_n35410,i_data[30]}),
    .sr(rst_pad),
    .q({open_n35416,\t/a/reg_writedat [30]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(C*~D)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111011111110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b31  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/a/MEM_aludat [31],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/a/MEM_aludat [31]}),
    .mi({open_n35428,i_data[31]}),
    .sr(rst_pad),
    .q({open_n35434,\t/a/reg_writedat [31]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(~C)"),
    //.LUT1("(~C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100001111),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \t/a/mem_wb/reg1_b1|t/a/mem_wb/reg1_b0  (
    .b({\t/a/MEM_op [1],open_n35437}),
    .c({\t/a/MEM_op [2],rst_pad}),
    .ce(\t/a/ex_mem/n0 ),
    .clk(clock_pad),
    .d({\t/a/MEM_op [0],open_n35438}),
    .mi(\t/a/MEM_op [1:0]),
    .f({_al_u251_o,\t/a/ex_mem/n0 }),
    .q(\t/a/WB_op [1:0]));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D"),
    //.LUTF1("0"),
    //.LUTG0("0"),
    //.LUTG1("~A*~B*~C*~D+~A*B*~C*~D"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011001100110011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \t/a/mem_wb/reg1_b2|t/a/mem_wb/reg1_b3  (
    .a({\t/a/WB_op [2],open_n35453}),
    .b({open_n35454,\t/a/MEM_op [4]}),
    .c({\t/a/WB_op [4],open_n35455}),
    .ce(\t/a/ex_mem/n0 ),
    .clk(clock_pad),
    .d({\t/a/WB_op [3],open_n35456}),
    .e({\t/a/WB_op [5],\t/a/MEM_op [3]}),
    .mi({\t/a/MEM_op [2],\t/a/MEM_op [3]}),
    .f({_al_u1793_o,_al_u252_o}),
    .q({\t/a/WB_op [2],\t/a/WB_op [3]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .MODE(),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \t/a/mem_wb/reg1_b4  (
    .ce(\t/a/ex_mem/n0 ),
    .clk(clock_pad),
    .mi({open_n35484,\t/a/MEM_op [4]}),
    .q({open_n35502,\t/a/WB_op [4]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("0"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("D*B*~C*~A+D*B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b1000010000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg2_b2|t/a/mem_wb/reg2_b0  (
    .a({\t/a/MEM_rd [2],_al_u1967_o}),
    .b({_al_u1969_o,\t/a/MEM_rd [0]}),
    .c({\t/a/EX_rs2 [2],\t/a/MEM_rd [1]}),
    .clk(clock_pad),
    .d({_al_u1968_o,\t/a/EX_rs2 [0]}),
    .e({_al_u1970_o,\t/a/EX_rs2 [1]}),
    .mi({\t/a/MEM_rd [2],\t/a/MEM_rd [0]}),
    .sr(rst_pad),
    .f({\t/a/n24_lutinv ,_al_u1968_o}),
    .q({\t/a/WB_rd [2],\t/a/WB_rd [0]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*((~0*B)*~(A)*~(D)+(~0*B)*A*~(D)+~((~0*B))*A*D+(~0*B)*A*D))"),
    //.LUT1("~(C*((~1*B)*~(A)*~(D)+(~1*B)*A*~(D)+~((~1*B))*A*D+(~1*B)*A*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101111100111111),
    .INIT_LUT1(16'b0101111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/regwritecs_reg  (
    .a({_al_u251_o,_al_u251_o}),
    .b({_al_u290_o,_al_u290_o}),
    .c({_al_u252_o,_al_u252_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_op [5],\t/a/MEM_op [5]}),
    .mi({open_n35530,\t/a/MEM_op [6]}),
    .sr(rst_pad),
    .q({open_n35536,\t/a/WB_regwritecs }));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1100110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b0|t/a/regfile/reg0_b9  (
    .a({open_n35537,\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/a/WB_regwritecs ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({open_n35538,\t/a/regfile/regfile$1$ [9]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/n46 [0],\t/a/regfile/regfile$0$ [9]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b0_sel_is_3_o ,_al_u1052_o}),
    .q({\t/a/regfile/regfile$0$ [0],\t/a/regfile/regfile$0$ [9]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*D*C*A*B)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*D*C*A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b1000|t/a/regfile/reg0_b999  (
    .a({\t/a/WB_rd [0],\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({_al_u256_o,\t/a/ID_rs2$1$_placeOpt_11 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2$2$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$30$ [7]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$31$ [7]}),
    .mi(\t/a/reg_writedat [8:7]),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b1000_sel_is_3_o ,_al_u1107_o}),
    .q(\t/a/regfile/regfile$31$ [8:7]));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000010101010),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0000000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b1001|t/a/regfile/reg0_b996  (
    .a({\t/a/reg_writedat [9],\t/a/ID_rs2$0$_placeOpt_10 }),
    .b({\t/a/MEM_aludat [9],\t/a/ID_rs2$1$_placeOpt_13 }),
    .c({open_n35567,\t/a/ID_rs2$2$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2614_o,\t/a/regfile/regfile$30$ [4]}),
    .e({_al_u2616_o_placeOpt_3,\t/a/regfile/regfile$31$ [4]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u2718_o,_al_u1170_o}),
    .q({\t/a/regfile/regfile$31$ [9],\t/a/regfile/regfile$31$ [4]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101010000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b1002|t/a/regfile/reg0_b995  (
    .a({_al_u2606_o_placeOpt_2,\t/a/ID_rs2$0$_placeOpt_16 }),
    .b({_al_u2610_o_placeOpt_2,\t/a/ID_rs2$1$_placeOpt_3 }),
    .c({\t/a/reg_writedat [10],\t/a/regfile/regfile$30$ [3]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [10],\t/a/regfile/regfile$31$ [3]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u2711_o,_al_u1177_o}),
    .q({\t/a/regfile/regfile$31$ [10],\t/a/regfile/regfile$31$ [3]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011000100100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b101|t/a/regfile/reg0_b99  (
    .a({_al_u2616_o,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({_al_u2614_o,\t/a/ID_rs2$1$_placeOpt_11 }),
    .c({\t/a/MEM_aludat [5],\t/a/regfile/regfile$2$ [3]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [5],\t/a/regfile/regfile$3$ [3]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u2740_o,_al_u1189_o}),
    .q({\t/a/regfile/regfile$3$ [5],\t/a/regfile/regfile$3$ [3]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b102|t/a/regfile/reg0_b98  (
    .a({_al_u2614_o,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({_al_u2616_o,\t/a/ID_rs2$1$_placeOpt_11 }),
    .c({\t/a/MEM_aludat [6],\t/a/regfile/regfile$2$ [2]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [6],\t/a/regfile/regfile$3$ [2]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u2733_o,_al_u1242_o}),
    .q({\t/a/regfile/regfile$3$ [6],\t/a/regfile/regfile$3$ [2]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0010001000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b103|t/a/regfile/reg0_b97  (
    .a({\t/a/MEM_aludat [7],\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({_al_u2614_o,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/reg_writedat [7],\t/a/regfile/regfile$2$ [1]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/regfile/regfile$3$ [1]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u2726_o,_al_u1473_o}),
    .q({\t/a/regfile/regfile$3$ [7],\t/a/regfile/regfile$3$ [1]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b107|t/a/regfile/reg0_b126  (
    .a({_al_u2606_o_placeOpt_3,_al_u2606_o_placeOpt_3}),
    .b({_al_u2610_o_placeOpt_3,_al_u2610_o_placeOpt_3}),
    .c({\t/a/MEM_aludat [11],\t/a/MEM_aludat [30]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [11],\t/a/reg_writedat [30]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u2703_o,_al_u2619_o}),
    .q({\t/a/regfile/regfile$3$ [11],\t/a/regfile/regfile$3$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b108|t/a/regfile/reg0_b125  (
    .a({_al_u2606_o_placeOpt_3,_al_u2606_o_placeOpt_3}),
    .b({_al_u2610_o_placeOpt_3,_al_u2610_o_placeOpt_3}),
    .c({\t/a/MEM_aludat [12],\t/a/MEM_aludat [29]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [12],\t/a/reg_writedat [29]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u2699_o,_al_u2623_o}),
    .q({\t/a/regfile/regfile$3$ [12],\t/a/regfile/regfile$3$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b109|t/a/regfile/reg0_b122  (
    .a({_al_u2606_o_placeOpt_3,_al_u2606_o_placeOpt_3}),
    .b({_al_u2610_o_placeOpt_3,_al_u2610_o_placeOpt_3}),
    .c({\t/a/MEM_aludat [13],\t/a/MEM_aludat [26]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [13],\t/a/reg_writedat [26]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u2695_o,_al_u2635_o}),
    .q({\t/a/regfile/regfile$3$ [13],\t/a/regfile/regfile$3$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b10|t/a/regfile/reg0_b8  (
    .a({_al_u2614_o_placeOpt_3,\t/a/ID_rs2$0$_placeOpt_3 }),
    .b({_al_u2616_o_placeOpt_3,\t/a/ID_rs2$1$_placeOpt_16 }),
    .c({\t/a/MEM_aludat [10],\t/a/regfile/regfile$1$ [8]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [10],\t/a/regfile/regfile$0$ [8]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u2714_o,_al_u1083_o}),
    .q({\t/a/regfile/regfile$0$ [10],\t/a/regfile/regfile$0$ [8]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101010000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b110|t/a/regfile/reg0_b121  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/reg_writedat [14],\t/a/MEM_aludat [25]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [14],\t/a/reg_writedat [25]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u2689_o,_al_u2639_o}),
    .q({\t/a/regfile/regfile$3$ [14],\t/a/regfile/regfile$3$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b111|t/a/regfile/reg0_b118  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/MEM_aludat [15],\t/a/MEM_aludat [22]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [15],\t/a/reg_writedat [22]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u2681_o,_al_u2651_o}),
    .q({\t/a/regfile/regfile$3$ [15],\t/a/regfile/regfile$3$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0100010101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b112|t/a/regfile/reg0_b117  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({\t/a/MEM_aludat [16],_al_u2610_o}),
    .c({_al_u2610_o,\t/a/MEM_aludat [21]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [16],\t/a/reg_writedat [21]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u2675_o,_al_u2655_o}),
    .q({\t/a/regfile/regfile$3$ [16],\t/a/regfile/regfile$3$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101010000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b113|t/a/regfile/reg0_b114  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/reg_writedat [17],\t/a/MEM_aludat [18]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [17],\t/a/reg_writedat [18]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u2671_o,_al_u2667_o}),
    .q({\t/a/regfile/regfile$3$ [17],\t/a/regfile/regfile$3$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b11|t/a/regfile/reg0_b7  (
    .a({_al_u2066_o,\t/a/ID_rs2$0$_placeOpt_14 }),
    .b({\t/a/alu_B_select [1],\t/a/ID_rs2$1$_placeOpt_19 }),
    .c({\t/a/aluin/n10_lutinv ,\t/a/regfile/regfile$1$ [7]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [11],\t/a/regfile/regfile$0$ [7]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b11/B9 ,_al_u1094_o}),
    .q({\t/a/regfile/regfile$0$ [11],\t/a/regfile/regfile$0$ [7]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(D*~A*~(~C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0101000100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b12|t/a/regfile/reg0_b6  (
    .a({_al_u2063_o,\t/a/ID_rs2$0$_placeOpt_9 }),
    .b({\t/a/alu_B_select [1],\t/a/ID_rs2$1$_placeOpt_18 }),
    .c({\t/a/reg_writedat [12],\t/a/regfile/regfile$1$ [6]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/n10_lutinv ,\t/a/regfile/regfile$0$ [6]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b12/B9 ,_al_u1115_o}),
    .q({\t/a/regfile/regfile$0$ [12],\t/a/regfile/regfile$0$ [6]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b137|t/a/regfile/reg0_b145  (
    .a({_al_u1979_o,_al_u2048_o}),
    .b({\t/a/alu_B_select [1],\t/a/alu_B_select [1]}),
    .c({\t/a/aluin/n10_lutinv ,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [9],\t/a/reg_writedat [17]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b9/B9 ,\t/a/aluin/sel1_b17/B9 }),
    .q({\t/a/regfile/regfile$4$ [9],\t/a/regfile/regfile$4$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(D*~A*~(~C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0101000100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b13|t/a/regfile/reg0_b5  (
    .a({_al_u2060_o,\t/a/ID_rs2$0$_placeOpt_10 }),
    .b({\t/a/alu_B_select [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/reg_writedat [13],\t/a/regfile/regfile$1$ [5]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/n10_lutinv ,\t/a/regfile/regfile$0$ [5]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b13/B9 ,_al_u1136_o}),
    .q({\t/a/regfile/regfile$0$ [13],\t/a/regfile/regfile$0$ [5]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(D*~A*~(~C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0101000100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b143|t/a/regfile/reg0_b144  (
    .a({_al_u2054_o,_al_u2051_o}),
    .b({\t/a/alu_B_select [1],\t/a/alu_B_select [1]}),
    .c({\t/a/reg_writedat [15],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/n10_lutinv ,\t/a/reg_writedat [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b15/B9 ,\t/a/aluin/sel1_b16/B9 }),
    .q({\t/a/regfile/regfile$4$ [15],\t/a/regfile/regfile$4$ [16]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(D*~A*~(~C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0101000100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b14|t/a/regfile/reg0_b4  (
    .a({_al_u2057_o,\t/a/ID_rs2$0$_placeOpt_3 }),
    .b({\t/a/alu_B_select [1],\t/a/ID_rs2$1$_placeOpt_13 }),
    .c({\t/a/reg_writedat [14],\t/a/regfile/regfile$1$ [4]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/n10_lutinv ,\t/a/regfile/regfile$0$ [4]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b14/B9 ,_al_u1157_o}),
    .q({\t/a/regfile/regfile$0$ [14],\t/a/regfile/regfile$0$ [4]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~A*~(~C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101000100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b15|t/a/regfile/reg0_b31  (
    .a({_al_u1877_o,\t/a/ID_rs1$0$_placeOpt_20 }),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1$1$_placeOpt_20 }),
    .c({\t/a/reg_writedat [15],\t/a/regfile/regfile$0$ [31]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$1$ [31]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b15/B0 ,_al_u493_o}),
    .q({\t/a/regfile/regfile$0$ [15],\t/a/regfile/regfile$0$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101010000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b162|t/a/regfile/reg0_b177  (
    .a({_al_u2606_o,\t/a/ID_rs1$0$_placeOpt_14 }),
    .b({_al_u2610_o,\t/a/ID_rs1$1$_placeOpt_14 }),
    .c({\t/a/reg_writedat [2],\t/a/regfile/regfile$4$ [17]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [2],\t/a/regfile/regfile$5$ [17]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u2754_o,_al_u817_o}),
    .q({\t/a/regfile/regfile$5$ [2],\t/a/regfile/regfile$5$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101010000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b163|t/a/regfile/reg0_b176  (
    .a({_al_u2606_o,\t/a/ID_rs1$0$_placeOpt_21 }),
    .b({_al_u2610_o,\t/a/ID_rs1$1$_placeOpt_21 }),
    .c({\t/a/reg_writedat [3],\t/a/regfile/regfile$4$ [16]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [3],\t/a/regfile/regfile$5$ [16]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u2749_o,_al_u848_o}),
    .q({\t/a/regfile/regfile$5$ [3],\t/a/regfile/regfile$5$ [16]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~A*~(~C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101000100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b16|t/a/regfile/reg0_b30  (
    .a({_al_u1874_o,\t/a/ID_rs1$0$_placeOpt_1 }),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1$1$_placeOpt_1 }),
    .c({\t/a/reg_writedat [16],\t/a/regfile/regfile$0$ [30]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$1$ [30]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b16/B0 ,_al_u504_o}),
    .q({\t/a/regfile/regfile$0$ [16],\t/a/regfile/regfile$0$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~A*~(~C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101000100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b17|t/a/regfile/reg0_b3  (
    .a({_al_u1871_o,\t/a/ID_rs1$0$_placeOpt_15 }),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1$1$_placeOpt_15 }),
    .c({\t/a/reg_writedat [17],\t/a/regfile/regfile$0$ [3]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$1$ [3]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b17/B0 ,_al_u462_o}),
    .q({\t/a/regfile/regfile$0$ [17],\t/a/regfile/regfile$0$ [3]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b18|t/a/regfile/reg0_b29  (
    .a({\t/a/ID_rs1$0$_placeOpt_21 ,\t/a/ID_rs1$0$_placeOpt_21 }),
    .b({\t/a/ID_rs1$1$_placeOpt_21 ,\t/a/ID_rs1$1$_placeOpt_21 }),
    .c({\t/a/regfile/regfile$0$ [18],\t/a/regfile/regfile$0$ [29]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [18],\t/a/regfile/regfile$1$ [29]}),
    .mi({\t/a/reg_writedat [18],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u808_o,_al_u556_o}),
    .q({\t/a/regfile/regfile$0$ [18],\t/a/regfile/regfile$0$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b193|t/a/regfile/reg0_b223  (
    .a({_al_u1895_o,\t/a/ID_rs1$0$_placeOpt_16 }),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1$1$_placeOpt_20 }),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [31]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [1],\t/a/regfile/regfile$7$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b1/B0 ,_al_u492_o}),
    .q({\t/a/regfile/regfile$6$ [1],\t/a/regfile/regfile$6$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b197|t/a/regfile/reg0_b222  (
    .a({_al_u1817_o,\t/a/ID_rs1$0$_placeOpt_20 }),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1$1$_placeOpt_20 }),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [30]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [5],\t/a/regfile/regfile$7$ [30]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b5/B0 ,_al_u503_o}),
    .q({\t/a/regfile/regfile$6$ [5],\t/a/regfile/regfile$6$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b198|t/a/regfile/reg0_b221  (
    .a({_al_u1814_o,\t/a/ID_rs1$0$_placeOpt_20 }),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1$1$_placeOpt_20 }),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [29]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [6],\t/a/regfile/regfile$7$ [29]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b6/B0 ,_al_u555_o}),
    .q({\t/a/regfile/regfile$6$ [6],\t/a/regfile/regfile$6$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~A*~(~C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b199|t/a/regfile/reg0_b220  (
    .a({_al_u1811_o,\t/a/ID_rs1$0$_placeOpt_20 }),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1$1$_placeOpt_20 }),
    .c({\t/a/reg_writedat [7],\t/a/regfile/regfile$6$ [28]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$7$ [28]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b7/B0 ,_al_u566_o}),
    .q({\t/a/regfile/regfile$6$ [7],\t/a/regfile/regfile$6$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b19|t/a/regfile/reg0_b28  (
    .a({\t/a/ID_rs1$0$_placeOpt_14 ,\t/a/ID_rs1$0$_placeOpt_14 }),
    .b({\t/a/ID_rs1$1$_placeOpt_14 ,\t/a/ID_rs1$1$_placeOpt_14 }),
    .c({\t/a/regfile/regfile$0$ [19],\t/a/regfile/regfile$0$ [28]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [19],\t/a/regfile/regfile$1$ [28]}),
    .mi({\t/a/reg_writedat [19],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u777_o,_al_u567_o}),
    .q({\t/a/regfile/regfile$0$ [19],\t/a/regfile/regfile$0$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0011000100100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b1|t/a/regfile/reg0_b27  (
    .a({_al_u2616_o,\t/a/ID_rs1$0$_placeOpt_16 }),
    .b({_al_u2614_o,\t/a/ID_rs1$1$_placeOpt_16 }),
    .c({\t/a/MEM_aludat [1],\t/a/regfile/regfile$0$ [27]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [1],\t/a/regfile/regfile$1$ [27]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u2764_o,_al_u598_o}),
    .q({\t/a/regfile/regfile$0$ [1],\t/a/regfile/regfile$0$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b200|t/a/regfile/reg0_b219  (
    .a({_al_u1808_o,\t/a/ID_rs1$0$_placeOpt_10 }),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [27]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [8],\t/a/regfile/regfile$7$ [27]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b8/B0 ,_al_u597_o}),
    .q({\t/a/regfile/regfile$6$ [8],\t/a/regfile/regfile$6$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b201|t/a/regfile/reg0_b218  (
    .a({\t/a/ID_rs1$0$_placeOpt_12 ,\t/a/ID_rs1$0$_placeOpt_12 }),
    .b({\t/a/ID_rs1$1$_placeOpt_12 ,\t/a/ID_rs1$1$_placeOpt_12 }),
    .c({\t/a/regfile/regfile$6$ [9],\t/a/regfile/regfile$6$ [26]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [9],\t/a/regfile/regfile$7$ [26]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u345_o,_al_u608_o}),
    .q({\t/a/regfile/regfile$6$ [9],\t/a/regfile/regfile$6$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b202|t/a/regfile/reg0_b217  (
    .a({\t/a/ID_rs1$0$_placeOpt_3 ,\t/a/ID_rs1$0$_placeOpt_3 }),
    .b({\t/a/ID_rs1$1$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$6$ [10],\t/a/regfile/regfile$6$ [25]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [10],\t/a/regfile/regfile$7$ [25]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u965_o,_al_u629_o}),
    .q({\t/a/regfile/regfile$6$ [10],\t/a/regfile/regfile$6$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b203|t/a/regfile/reg0_b216  (
    .a({\t/a/ID_rs1$0$_placeOpt_14 ,\t/a/ID_rs1$0$_placeOpt_14 }),
    .b({\t/a/ID_rs1$1$_placeOpt_14 ,\t/a/ID_rs1$1$_placeOpt_14 }),
    .c({\t/a/regfile/regfile$7$ [11],\t/a/regfile/regfile$6$ [24]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$6$ [11],\t/a/regfile/regfile$7$ [24]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u954_o,_al_u650_o}),
    .q({\t/a/regfile/regfile$6$ [11],\t/a/regfile/regfile$6$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b204|t/a/regfile/reg0_b215  (
    .a({\t/a/ID_rs1$0$_placeOpt_9 ,\t/a/ID_rs1$0$_placeOpt_9 }),
    .b({\t/a/ID_rs1$1$_placeOpt_9 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .c({\t/a/regfile/regfile$6$ [12],\t/a/regfile/regfile$6$ [23]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [12],\t/a/regfile/regfile$7$ [23]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u923_o,_al_u671_o}),
    .q({\t/a/regfile/regfile$6$ [12],\t/a/regfile/regfile$6$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b205|t/a/regfile/reg0_b214  (
    .a({\t/a/ID_rs1$0$_placeOpt_3 ,\t/a/ID_rs1$0$_placeOpt_3 }),
    .b({\t/a/ID_rs1$1$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$6$ [13],\t/a/regfile/regfile$6$ [22]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [13],\t/a/regfile/regfile$7$ [22]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u912_o,_al_u702_o}),
    .q({\t/a/regfile/regfile$6$ [13],\t/a/regfile/regfile$6$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b206|t/a/regfile/reg0_b213  (
    .a({\t/a/ID_rs1$0$_placeOpt_11 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .b({\t/a/ID_rs1$1$_placeOpt_11 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$6$ [14],\t/a/regfile/regfile$6$ [21]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [14],\t/a/regfile/regfile$7$ [21]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u881_o,_al_u713_o}),
    .q({\t/a/regfile/regfile$6$ [14],\t/a/regfile/regfile$6$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b207|t/a/regfile/reg0_b212  (
    .a({\t/a/ID_rs1$0$_placeOpt_17 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .b({\t/a/ID_rs1$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$7$ [15],\t/a/regfile/regfile$6$ [20]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$6$ [15],\t/a/regfile/regfile$7$ [20]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u860_o,_al_u744_o}),
    .q({\t/a/regfile/regfile$6$ [15],\t/a/regfile/regfile$6$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b208|t/a/regfile/reg0_b211  (
    .a({\t/a/ID_rs1$0$_placeOpt_17 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .b({\t/a/ID_rs1$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$6$ [16],\t/a/regfile/regfile$6$ [19]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [16],\t/a/regfile/regfile$7$ [19]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u849_o,_al_u776_o}),
    .q({\t/a/regfile/regfile$6$ [16],\t/a/regfile/regfile$6$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b209|t/a/regfile/reg0_b210  (
    .a({\t/a/ID_rs1$0$_placeOpt_17 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .b({\t/a/ID_rs1$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$6$ [17],\t/a/regfile/regfile$6$ [18]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [17],\t/a/regfile/regfile$7$ [18]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u818_o,_al_u807_o}),
    .q({\t/a/regfile/regfile$6$ [17],\t/a/regfile/regfile$6$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b20|t/a/regfile/reg0_b26  (
    .a({\t/a/ID_rs1$0$_placeOpt_9 ,\t/a/ID_rs1$0$_placeOpt_9 }),
    .b({\t/a/ID_rs1$1$_placeOpt_9 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .c({\t/a/regfile/regfile$0$ [20],\t/a/regfile/regfile$0$ [26]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [20],\t/a/regfile/regfile$1$ [26]}),
    .mi({\t/a/reg_writedat [20],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u745_o,_al_u609_o}),
    .q({\t/a/regfile/regfile$0$ [20],\t/a/regfile/regfile$0$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b21|t/a/regfile/reg0_b25  (
    .a({\t/a/ID_rs1$0$_placeOpt_14 ,\t/a/ID_rs1$0$_placeOpt_14 }),
    .b({\t/a/ID_rs1$1$_placeOpt_14 ,\t/a/ID_rs1$1$_placeOpt_14 }),
    .c({\t/a/regfile/regfile$0$ [21],\t/a/regfile/regfile$0$ [25]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [21],\t/a/regfile/regfile$1$ [25]}),
    .mi({\t/a/reg_writedat [21],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u714_o,_al_u630_o}),
    .q({\t/a/regfile/regfile$0$ [21],\t/a/regfile/regfile$0$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b225|t/a/regfile/reg0_b255  (
    .a({\t/a/regfile/regfile$6$ [1],\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/a/regfile/regfile$7$ [1],\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/regfile/regfile$6$ [31]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/regfile/regfile$7$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u755_o,_al_u1198_o}),
    .q({\t/a/regfile/regfile$7$ [1],\t/a/regfile/regfile$7$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b226|t/a/regfile/reg0_b254  (
    .a({\t/a/regfile/regfile$7$ [2],\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/a/regfile/regfile$6$ [2],\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/regfile/regfile$6$ [30]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/regfile/regfile$7$ [30]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u524_o,_al_u1229_o}),
    .q({\t/a/regfile/regfile$7$ [2],\t/a/regfile/regfile$7$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b227|t/a/regfile/reg0_b253  (
    .a({_al_u1829_o,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs2$1$_placeOpt_11 }),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [29]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [3],\t/a/regfile/regfile$7$ [29]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b3/B0 ,_al_u1261_o}),
    .q({\t/a/regfile/regfile$7$ [3],\t/a/regfile/regfile$7$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b228|t/a/regfile/reg0_b252  (
    .a({_al_u1820_o,\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [28]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [4],\t/a/regfile/regfile$7$ [28]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b4/B0 ,_al_u1292_o}),
    .q({\t/a/regfile/regfile$7$ [4],\t/a/regfile/regfile$7$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b229|t/a/regfile/reg0_b251  (
    .a({\t/a/regfile/regfile$7$ [5],\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/regfile/regfile$6$ [5],\t/a/ID_rs2$1$_placeOpt_11 }),
    .c({\t/a/ID_rs1$1$_placeOpt_10 ,\t/a/regfile/regfile$6$ [27]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_10 ,\t/a/regfile/regfile$7$ [27]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u419_o,_al_u1303_o}),
    .q({\t/a/regfile/regfile$7$ [5],\t/a/regfile/regfile$7$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b22|t/a/regfile/reg0_b24  (
    .a({\t/a/ID_rs1$0$_placeOpt_3 ,\t/a/ID_rs1$0$_placeOpt_3 }),
    .b({\t/a/ID_rs1$1$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$0$ [22],\t/a/regfile/regfile$0$ [24]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [22],\t/a/regfile/regfile$1$ [24]}),
    .mi({\t/a/reg_writedat [22],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u703_o,_al_u651_o}),
    .q({\t/a/regfile/regfile$0$ [22],\t/a/regfile/regfile$0$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b230|t/a/regfile/reg0_b250  (
    .a({\t/a/ID_rs1$0$_placeOpt_12 ,\t/a/ID_rs2$0$_placeOpt_11 }),
    .b({\t/a/ID_rs1$1$_placeOpt_12 ,\t/a/ID_rs2$1$_placeOpt_9 }),
    .c({\t/a/regfile/regfile$6$ [6],\t/a/regfile/regfile$6$ [26]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [6],\t/a/regfile/regfile$7$ [26]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u398_o,_al_u1334_o}),
    .q({\t/a/regfile/regfile$7$ [6],\t/a/regfile/regfile$7$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b231|t/a/regfile/reg0_b249  (
    .a({\t/a/regfile/regfile$6$ [7],\t/a/ID_rs2$0$_placeOpt_16 }),
    .b({\t/a/regfile/regfile$7$ [7],\t/a/ID_rs2$1$_placeOpt_3 }),
    .c({\t/a/ID_rs1$0$_placeOpt_2 ,\t/a/regfile/regfile$6$ [25]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_2 ,\t/a/regfile/regfile$7$ [25]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u387_o,_al_u1345_o}),
    .q({\t/a/regfile/regfile$7$ [7],\t/a/regfile/regfile$7$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b232|t/a/regfile/reg0_b248  (
    .a({\t/a/regfile/regfile$6$ [8],\t/a/ID_rs2$0$_placeOpt_14 }),
    .b({\t/a/regfile/regfile$7$ [8],\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/ID_rs1$0$_placeOpt_3 ,\t/a/regfile/regfile$6$ [24]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_3 ,\t/a/regfile/regfile$7$ [24]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u356_o,_al_u1366_o}),
    .q({\t/a/regfile/regfile$7$ [8],\t/a/regfile/regfile$7$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b233|t/a/regfile/reg0_b247  (
    .a({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs2$0$_placeOpt_20 }),
    .b({\t/a/ID_rs2$1$_placeOpt_21 ,\t/a/ID_rs2$1$_placeOpt_21 }),
    .c({\t/a/regfile/regfile$7$ [9],\t/a/regfile/regfile$6$ [23]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$6$ [9],\t/a/regfile/regfile$7$ [23]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1051_o,_al_u1397_o}),
    .q({\t/a/regfile/regfile$7$ [9],\t/a/regfile/regfile$7$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b234|t/a/regfile/reg0_b246  (
    .a({\t/a/ID_rs2$0$_placeOpt_8 ,\t/a/ID_rs2$0$_placeOpt_8 }),
    .b({\t/a/ID_rs2$1$_placeOpt_16 ,\t/a/ID_rs2$1$_placeOpt_16 }),
    .c({\t/a/regfile/regfile$7$ [10],\t/a/regfile/regfile$6$ [22]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$6$ [10],\t/a/regfile/regfile$7$ [22]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1691_o,_al_u1408_o}),
    .q({\t/a/regfile/regfile$7$ [10],\t/a/regfile/regfile$7$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b235|t/a/regfile/reg0_b245  (
    .a({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs2$0$_placeOpt_12 }),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_5 }),
    .c({\t/a/regfile/regfile$6$ [11],\t/a/regfile/regfile$6$ [21]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [11],\t/a/regfile/regfile$7$ [21]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1660_o,_al_u1439_o}),
    .q({\t/a/regfile/regfile$7$ [11],\t/a/regfile/regfile$7$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b236|t/a/regfile/reg0_b244  (
    .a({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs2$0$_placeOpt_20 }),
    .b({\t/a/ID_rs2$1$_placeOpt_10 ,\t/a/ID_rs2$1$_placeOpt_10 }),
    .c({\t/a/regfile/regfile$6$ [12],\t/a/regfile/regfile$6$ [20]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [12],\t/a/regfile/regfile$7$ [20]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1649_o,_al_u1450_o}),
    .q({\t/a/regfile/regfile$7$ [12],\t/a/regfile/regfile$7$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b237|t/a/regfile/reg0_b243  (
    .a({\t/a/ID_rs2$0$_placeOpt_19 ,\t/a/ID_rs2$0$_placeOpt_19 }),
    .b({\t/a/ID_rs2$1$_placeOpt_14 ,\t/a/ID_rs2$1$_placeOpt_14 }),
    .c({\t/a/regfile/regfile$7$ [13],\t/a/regfile/regfile$6$ [19]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$6$ [13],\t/a/regfile/regfile$7$ [19]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1618_o,_al_u1492_o}),
    .q({\t/a/regfile/regfile$7$ [13],\t/a/regfile/regfile$7$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b238|t/a/regfile/reg0_b242  (
    .a({\t/a/ID_rs2$0$_placeOpt_13 ,\t/a/ID_rs2$0$_placeOpt_13 }),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs2$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$7$ [14],\t/a/regfile/regfile$6$ [18]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$6$ [14],\t/a/regfile/regfile$7$ [18]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1597_o,_al_u1513_o}),
    .q({\t/a/regfile/regfile$7$ [14],\t/a/regfile/regfile$7$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b239|t/a/regfile/reg0_b241  (
    .a({\t/a/ID_rs2$0$_placeOpt_13 ,\t/a/ID_rs2$0$_placeOpt_13 }),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs2$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$6$ [15],\t/a/regfile/regfile$6$ [17]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [15],\t/a/regfile/regfile$7$ [17]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1586_o,_al_u1544_o}),
    .q({\t/a/regfile/regfile$7$ [15],\t/a/regfile/regfile$7$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b256|t/a/regfile/reg0_b287  (
    .a({_al_u254_o,_al_u498_o}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1$0$_placeOpt_16 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1$1$_placeOpt_16 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$8$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$9$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b256_sel_is_3_o ,_al_u499_o}),
    .q({\t/a/regfile/regfile$8$ [0],\t/a/regfile/regfile$8$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b257|t/a/regfile/reg0_b286  (
    .a({_al_u761_o,_al_u509_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/ID_rs1$0$_placeOpt_16 }),
    .c({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/ID_rs1$1$_placeOpt_16 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [1],\t/a/regfile/regfile$8$ [30]}),
    .e({\t/a/regfile/regfile$9$ [1],\t/a/regfile/regfile$9$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u762_o,_al_u510_o}),
    .q({\t/a/regfile/regfile$8$ [1],\t/a/regfile/regfile$8$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b258|t/a/regfile/reg0_b285  (
    .a({_al_u530_o,_al_u561_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_12 ,\t/a/ID_rs1$0$_placeOpt_12 }),
    .c({\t/a/ID_rs1$1$_placeOpt_12 ,\t/a/ID_rs1$1$_placeOpt_12 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [2],\t/a/regfile/regfile$8$ [29]}),
    .e({\t/a/regfile/regfile$9$ [2],\t/a/regfile/regfile$9$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u531_o,_al_u562_o}),
    .q({\t/a/regfile/regfile$8$ [2],\t/a/regfile/regfile$8$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b259|t/a/regfile/reg0_b284  (
    .a({_al_u467_o,_al_u572_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_13 }),
    .c({\t/a/regfile/regfile$8$ [3],\t/a/ID_rs1$1$_placeOpt_13 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/regfile/regfile$8$ [28]}),
    .e({\t/a/regfile/regfile$9$ [3],\t/a/regfile/regfile$9$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u468_o,_al_u573_o}),
    .q({\t/a/regfile/regfile$8$ [3],\t/a/regfile/regfile$8$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b260|t/a/regfile/reg0_b283  (
    .a({_al_u456_o,_al_u603_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_13 }),
    .c({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/ID_rs1$1$_placeOpt_13 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [4],\t/a/regfile/regfile$8$ [27]}),
    .e({\t/a/regfile/regfile$9$ [4],\t/a/regfile/regfile$9$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u457_o,_al_u604_o}),
    .q({\t/a/regfile/regfile$8$ [4],\t/a/regfile/regfile$8$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b261|t/a/regfile/reg0_b282  (
    .a({_al_u425_o,_al_u614_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_9 ,\t/a/ID_rs1$0$_placeOpt_9 }),
    .c({\t/a/ID_rs1$1$_placeOpt_9 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [5],\t/a/regfile/regfile$8$ [26]}),
    .e({\t/a/regfile/regfile$9$ [5],\t/a/regfile/regfile$9$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u426_o,_al_u615_o}),
    .q({\t/a/regfile/regfile$8$ [5],\t/a/regfile/regfile$8$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b262|t/a/regfile/reg0_b281  (
    .a({_al_u404_o,_al_u635_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_17 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$8$ [6],\t/a/ID_rs1$1$_placeOpt_17 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_17 ,\t/a/regfile/regfile$8$ [25]}),
    .e({\t/a/regfile/regfile$9$ [6],\t/a/regfile/regfile$9$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u405_o,_al_u636_o}),
    .q({\t/a/regfile/regfile$8$ [6],\t/a/regfile/regfile$8$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b263|t/a/regfile/reg0_b280  (
    .a({_al_u393_o,_al_u656_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_19 ,\t/a/ID_rs1$0$_placeOpt_19 }),
    .c({\t/a/ID_rs1$1$_placeOpt_19 ,\t/a/ID_rs1$1$_placeOpt_19 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [7],\t/a/regfile/regfile$8$ [24]}),
    .e({\t/a/regfile/regfile$9$ [7],\t/a/regfile/regfile$9$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u394_o,_al_u657_o}),
    .q({\t/a/regfile/regfile$8$ [7],\t/a/regfile/regfile$8$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b264|t/a/regfile/reg0_b279  (
    .a({_al_u362_o,_al_u677_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_12 ,\t/a/ID_rs1$0$_placeOpt_12 }),
    .c({\t/a/ID_rs1$1$_placeOpt_12 ,\t/a/ID_rs1$1$_placeOpt_12 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [8],\t/a/regfile/regfile$8$ [23]}),
    .e({\t/a/regfile/regfile$9$ [8],\t/a/regfile/regfile$9$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u363_o,_al_u678_o}),
    .q({\t/a/regfile/regfile$8$ [8],\t/a/regfile/regfile$8$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b265|t/a/regfile/reg0_b278  (
    .a({_al_u351_o,_al_u708_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_13 }),
    .c({\t/a/regfile/regfile$8$ [9],\t/a/ID_rs1$1$_placeOpt_13 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/regfile/regfile$8$ [22]}),
    .e({\t/a/regfile/regfile$9$ [9],\t/a/regfile/regfile$9$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u352_o,_al_u709_o}),
    .q({\t/a/regfile/regfile$8$ [9],\t/a/regfile/regfile$8$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b266|t/a/regfile/reg0_b277  (
    .a({_al_u971_o,_al_u719_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .c({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/ID_rs1$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [10],\t/a/regfile/regfile$8$ [21]}),
    .e({\t/a/regfile/regfile$9$ [10],\t/a/regfile/regfile$9$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u972_o,_al_u720_o}),
    .q({\t/a/regfile/regfile$8$ [10],\t/a/regfile/regfile$8$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b267|t/a/regfile/reg0_b276  (
    .a({_al_u960_o,_al_u750_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_17 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .c({\t/a/ID_rs1$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [11],\t/a/regfile/regfile$8$ [20]}),
    .e({\t/a/regfile/regfile$9$ [11],\t/a/regfile/regfile$9$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u961_o,_al_u751_o}),
    .q({\t/a/regfile/regfile$8$ [11],\t/a/regfile/regfile$8$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b268|t/a/regfile/reg0_b275  (
    .a({_al_u929_o,_al_u782_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_17 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .c({\t/a/ID_rs1$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [12],\t/a/regfile/regfile$8$ [19]}),
    .e({\t/a/regfile/regfile$9$ [12],\t/a/regfile/regfile$9$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u930_o,_al_u783_o}),
    .q({\t/a/regfile/regfile$8$ [12],\t/a/regfile/regfile$8$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b269|t/a/regfile/reg0_b274  (
    .a({_al_u918_o,_al_u813_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_11 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .c({\t/a/ID_rs1$1$_placeOpt_11 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [13],\t/a/regfile/regfile$8$ [18]}),
    .e({\t/a/regfile/regfile$9$ [13],\t/a/regfile/regfile$9$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u919_o,_al_u814_o}),
    .q({\t/a/regfile/regfile$8$ [13],\t/a/regfile/regfile$8$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b270|t/a/regfile/reg0_b273  (
    .a({_al_u887_o,_al_u824_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_11 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .c({\t/a/ID_rs1$1$_placeOpt_11 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [14],\t/a/regfile/regfile$8$ [17]}),
    .e({\t/a/regfile/regfile$9$ [14],\t/a/regfile/regfile$9$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u888_o,_al_u825_o}),
    .q({\t/a/regfile/regfile$8$ [14],\t/a/regfile/regfile$8$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b271|t/a/regfile/reg0_b272  (
    .a({_al_u866_o,_al_u855_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_9 ,\t/a/ID_rs1$0$_placeOpt_9 }),
    .c({\t/a/ID_rs1$1$_placeOpt_9 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [15],\t/a/regfile/regfile$8$ [16]}),
    .e({\t/a/regfile/regfile$9$ [15],\t/a/regfile/regfile$9$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u867_o,_al_u856_o}),
    .q({\t/a/regfile/regfile$8$ [15],\t/a/regfile/regfile$8$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*~D*~C*A*B)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*~D*~C*A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b288|t/a/regfile/reg0_b319  (
    .a({\t/a/WB_rd [0],_al_u1204_o}),
    .b({_al_u254_o,\t/a/ID_rs2$0$_placeOpt_21 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2$1$_placeOpt_15 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$8$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$9$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b288_sel_is_3_o ,_al_u1205_o}),
    .q({\t/a/regfile/regfile$9$ [0],\t/a/regfile/regfile$9$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b289|t/a/regfile/reg0_b318  (
    .a({_al_u1477_o,_al_u1235_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/ID_rs2$0$_placeOpt_21 }),
    .c({\t/a/regfile/regfile$8$ [1],\t/a/ID_rs2$1$_placeOpt_15 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/regfile/regfile$8$ [30]}),
    .e({\t/a/regfile/regfile$9$ [1],\t/a/regfile/regfile$9$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1478_o,_al_u1236_o}),
    .q({\t/a/regfile/regfile$9$ [1],\t/a/regfile/regfile$9$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~B*~(C*~(0)*~(D)+C*0*~(D)+~(C)*0*D+C*0*D)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~B*~(C*~(1)*~(D)+C*1*~(D)+~(C)*1*D+C*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1000100010101000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b290|t/a/regfile/reg0_b317  (
    .a({_al_u1246_o,_al_u1267_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_9 ,\t/a/ID_rs2$0$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$8$ [2],\t/a/ID_rs2$1$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_11 ,\t/a/regfile/regfile$8$ [29]}),
    .e({\t/a/regfile/regfile$9$ [2],\t/a/regfile/regfile$9$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1247_o,_al_u1268_o}),
    .q({\t/a/regfile/regfile$9$ [2],\t/a/regfile/regfile$9$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1000101010001000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b291|t/a/regfile/reg0_b316  (
    .a({_al_u1193_o,_al_u1298_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_20 ,\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [0],\t/a/ID_rs2$1$_placeOpt_20 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [3],\t/a/regfile/regfile$8$ [28]}),
    .e({\t/a/regfile/regfile$9$ [3],\t/a/regfile/regfile$9$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1194_o,_al_u1299_o}),
    .q({\t/a/regfile/regfile$9$ [3],\t/a/regfile/regfile$9$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b292|t/a/regfile/reg0_b315  (
    .a({_al_u1162_o,_al_u1309_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/ID_rs2$0$_placeOpt_22 }),
    .c({\t/a/ID_rs2$1$_placeOpt_12 ,\t/a/ID_rs2$1$_placeOpt_12 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [4],\t/a/regfile/regfile$8$ [27]}),
    .e({\t/a/regfile/regfile$9$ [4],\t/a/regfile/regfile$9$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1163_o,_al_u1310_o}),
    .q({\t/a/regfile/regfile$9$ [4],\t/a/regfile/regfile$9$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b293|t/a/regfile/reg0_b314  (
    .a({_al_u1141_o,_al_u1340_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs2$0$_placeOpt_20 }),
    .c({\t/a/ID_rs2$1$_placeOpt_21 ,\t/a/ID_rs2$1$_placeOpt_21 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [5],\t/a/regfile/regfile$8$ [26]}),
    .e({\t/a/regfile/regfile$9$ [5],\t/a/regfile/regfile$9$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1142_o,_al_u1341_o}),
    .q({\t/a/regfile/regfile$9$ [5],\t/a/regfile/regfile$9$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b294|t/a/regfile/reg0_b313  (
    .a({_al_u1120_o,_al_u1351_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_17 ,\t/a/ID_rs2$0$_placeOpt_17 }),
    .c({\t/a/ID_rs2$1$_placeOpt_8 ,\t/a/ID_rs2$1$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [6],\t/a/regfile/regfile$8$ [25]}),
    .e({\t/a/regfile/regfile$9$ [6],\t/a/regfile/regfile$9$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1121_o,_al_u1352_o}),
    .q({\t/a/regfile/regfile$9$ [6],\t/a/regfile/regfile$9$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(D*~(~A*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(D*~(~A*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1011101000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1111111000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b295|t/a/regfile/reg0_b312  (
    .a({\t/a/ID_rs2$1$_placeOpt_20 ,_al_u1372_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/regfile/regfile$8$ [7],\t/a/ID_rs2$1$_placeOpt_20 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u1099_o,\t/a/regfile/regfile$8$ [24]}),
    .e({\t/a/regfile/regfile$9$ [7],\t/a/regfile/regfile$9$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1100_o,_al_u1373_o}),
    .q({\t/a/regfile/regfile$9$ [7],\t/a/regfile/regfile$9$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1000101010001000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b296|t/a/regfile/reg0_b311  (
    .a({_al_u1088_o,_al_u1403_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_9 ,\t/a/ID_rs2$0$_placeOpt_11 }),
    .c({\t/a/ID_rs2$0$_placeOpt_11 ,\t/a/ID_rs2$1$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [8],\t/a/regfile/regfile$8$ [23]}),
    .e({\t/a/regfile/regfile$9$ [8],\t/a/regfile/regfile$9$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1089_o,_al_u1404_o}),
    .q({\t/a/regfile/regfile$9$ [8],\t/a/regfile/regfile$9$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1000101010001000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b297|t/a/regfile/reg0_b310  (
    .a({_al_u1057_o,_al_u1414_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_20 ,\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [0],\t/a/ID_rs2$1$_placeOpt_20 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [9],\t/a/regfile/regfile$8$ [22]}),
    .e({\t/a/regfile/regfile$9$ [9],\t/a/regfile/regfile$9$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1058_o,_al_u1415_o}),
    .q({\t/a/regfile/regfile$9$ [9],\t/a/regfile/regfile$9$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b298|t/a/regfile/reg0_b309  (
    .a({_al_u1697_o,_al_u1445_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs2$0$_placeOpt_12 }),
    .c({\t/a/regfile/regfile$8$ [10],\t/a/ID_rs2$1$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/regfile/regfile$8$ [21]}),
    .e({\t/a/regfile/regfile$9$ [10],\t/a/regfile/regfile$9$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1698_o,_al_u1446_o}),
    .q({\t/a/regfile/regfile$9$ [10],\t/a/regfile/regfile$9$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b299|t/a/regfile/reg0_b308  (
    .a({_al_u1666_o,_al_u1456_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_13 ,\t/a/ID_rs2$0$_placeOpt_13 }),
    .c({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs2$1$_placeOpt_17 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [11],\t/a/regfile/regfile$8$ [20]}),
    .e({\t/a/regfile/regfile$9$ [11],\t/a/regfile/regfile$9$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1667_o,_al_u1457_o}),
    .q({\t/a/regfile/regfile$9$ [11],\t/a/regfile/regfile$9$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b2|t/a/regfile/reg0_b23  (
    .a({_al_u1862_o,\t/a/ID_rs1$0$_placeOpt_16 }),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$0$ [23]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [2],\t/a/regfile/regfile$1$ [23]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b2/B0 ,_al_u672_o}),
    .q({\t/a/regfile/regfile$0$ [2],\t/a/regfile/regfile$0$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b300|t/a/regfile/reg0_b307  (
    .a({_al_u1655_o,_al_u1498_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs2$0$_placeOpt_20 }),
    .c({\t/a/ID_rs2$1$_placeOpt_10 ,\t/a/ID_rs2$1$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [12],\t/a/regfile/regfile$8$ [19]}),
    .e({\t/a/regfile/regfile$9$ [12],\t/a/regfile/regfile$9$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1656_o,_al_u1499_o}),
    .q({\t/a/regfile/regfile$9$ [12],\t/a/regfile/regfile$9$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(B*~(~D*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(B*~(~D*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1100110001000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100110011001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b301|t/a/regfile/reg0_b306  (
    .a({\t/a/ID_rs2$0$_placeOpt_17 ,_al_u1519_o}),
    .b({_al_u1624_o,\t/a/ID_rs2$0$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$8$ [13],\t/a/ID_rs2$1$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_8 ,\t/a/regfile/regfile$8$ [18]}),
    .e({\t/a/regfile/regfile$9$ [13],\t/a/regfile/regfile$9$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1625_o,_al_u1520_o}),
    .q({\t/a/regfile/regfile$9$ [13],\t/a/regfile/regfile$9$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b302|t/a/regfile/reg0_b305  (
    .a({_al_u1603_o,_al_u1550_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_17 ,\t/a/ID_rs2$0$_placeOpt_17 }),
    .c({\t/a/ID_rs2$1$_placeOpt_8 ,\t/a/ID_rs2$1$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [14],\t/a/regfile/regfile$8$ [17]}),
    .e({\t/a/regfile/regfile$9$ [14],\t/a/regfile/regfile$9$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1604_o,_al_u1551_o}),
    .q({\t/a/regfile/regfile$9$ [14],\t/a/regfile/regfile$9$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b303|t/a/regfile/reg0_b304  (
    .a({_al_u1592_o,_al_u1561_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs2$0$_placeOpt_20 }),
    .c({\t/a/ID_rs2$1$_placeOpt_10 ,\t/a/ID_rs2$1$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [15],\t/a/regfile/regfile$8$ [16]}),
    .e({\t/a/regfile/regfile$9$ [15],\t/a/regfile/regfile$9$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1593_o,_al_u1562_o}),
    .q({\t/a/regfile/regfile$9$ [15],\t/a/regfile/regfile$9$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*~D*C*~B*A)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*~D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b320|t/a/regfile/reg0_b351  (
    .a({_al_u254_o,\t/a/ID_rs1$0$_placeOpt_16 }),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$10$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$11$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b320_sel_is_3_o ,_al_u498_o}),
    .q({\t/a/regfile/regfile$10$ [0],\t/a/regfile/regfile$10$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b321|t/a/regfile/reg0_b350  (
    .a({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/ID_rs1$0$_placeOpt_16 }),
    .b({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/ID_rs1$1$_placeOpt_16 }),
    .c({\t/a/ID_rs1$2$_placeOpt_6 ,\t/a/ID_rs1$2$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [1],\t/a/regfile/regfile$10$ [30]}),
    .e({\t/a/regfile/regfile$11$ [1],\t/a/regfile/regfile$11$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u761_o,_al_u509_o}),
    .q({\t/a/regfile/regfile$10$ [1],\t/a/regfile/regfile$10$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b322|t/a/regfile/reg0_b349  (
    .a({\t/a/ID_rs1$0$_placeOpt_12 ,\t/a/ID_rs1$0$_placeOpt_12 }),
    .b({\t/a/ID_rs1$1$_placeOpt_12 ,\t/a/ID_rs1$1$_placeOpt_12 }),
    .c({\t/a/ID_rs1$2$_placeOpt_8 ,\t/a/ID_rs1$2$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [2],\t/a/regfile/regfile$10$ [29]}),
    .e({\t/a/regfile/regfile$11$ [2],\t/a/regfile/regfile$11$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u530_o,_al_u561_o}),
    .q({\t/a/regfile/regfile$10$ [2],\t/a/regfile/regfile$10$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b323|t/a/regfile/reg0_b348  (
    .a({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_13 }),
    .b({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/ID_rs1$1$_placeOpt_13 }),
    .c({\t/a/ID_rs1$2$_placeOpt_4 ,\t/a/ID_rs1$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [3],\t/a/regfile/regfile$10$ [28]}),
    .e({\t/a/regfile/regfile$11$ [3],\t/a/regfile/regfile$11$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u467_o,_al_u572_o}),
    .q({\t/a/regfile/regfile$10$ [3],\t/a/regfile/regfile$10$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b324|t/a/regfile/reg0_b347  (
    .a({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_13 }),
    .b({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/ID_rs1$1$_placeOpt_13 }),
    .c({\t/a/ID_rs1$2$_placeOpt_4 ,\t/a/ID_rs1$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [4],\t/a/regfile/regfile$10$ [27]}),
    .e({\t/a/regfile/regfile$11$ [4],\t/a/regfile/regfile$11$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u456_o,_al_u603_o}),
    .q({\t/a/regfile/regfile$10$ [4],\t/a/regfile/regfile$10$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000011111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b325|t/a/regfile/reg0_b346  (
    .a({\t/a/ID_rs1$0$_placeOpt_9 ,\t/a/ID_rs1$0$_placeOpt_9 }),
    .b({\t/a/ID_rs1$1$_placeOpt_9 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .c({\t/a/regfile/regfile$10$ [5],\t/a/ID_rs1$2$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$2$_placeOpt_8 ,\t/a/regfile/regfile$10$ [26]}),
    .e({\t/a/regfile/regfile$11$ [5],\t/a/regfile/regfile$11$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u425_o,_al_u614_o}),
    .q({\t/a/regfile/regfile$10$ [5],\t/a/regfile/regfile$10$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b326|t/a/regfile/reg0_b345  (
    .a({\t/a/ID_rs1$0$_placeOpt_11 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .b({\t/a/ID_rs1$1$_placeOpt_11 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/ID_rs1$2$_placeOpt_5 ,\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [6],\t/a/regfile/regfile$10$ [25]}),
    .e({\t/a/regfile/regfile$11$ [6],\t/a/regfile/regfile$11$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u404_o,_al_u635_o}),
    .q({\t/a/regfile/regfile$10$ [6],\t/a/regfile/regfile$10$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~A*~(B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~A*~(B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0001010100010001),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0101010101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b327|t/a/regfile/reg0_b344  (
    .a({\t/a/ID_rs1 [2],\t/a/ID_rs1$0$_placeOpt_19 }),
    .b({\t/a/ID_rs1$1$_placeOpt_19 ,\t/a/ID_rs1$1$_placeOpt_19 }),
    .c({\t/a/ID_rs1$0$_placeOpt_19 ,\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [7],\t/a/regfile/regfile$10$ [24]}),
    .e({\t/a/regfile/regfile$11$ [7],\t/a/regfile/regfile$11$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u393_o,_al_u656_o}),
    .q({\t/a/regfile/regfile$10$ [7],\t/a/regfile/regfile$10$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b328|t/a/regfile/reg0_b343  (
    .a({\t/a/ID_rs1$0$_placeOpt_12 ,\t/a/ID_rs1$0$_placeOpt_12 }),
    .b({\t/a/ID_rs1$1$_placeOpt_12 ,\t/a/ID_rs1$1$_placeOpt_12 }),
    .c({\t/a/ID_rs1$2$_placeOpt_8 ,\t/a/ID_rs1$2$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [8],\t/a/regfile/regfile$10$ [23]}),
    .e({\t/a/regfile/regfile$11$ [8],\t/a/regfile/regfile$11$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u362_o,_al_u677_o}),
    .q({\t/a/regfile/regfile$10$ [8],\t/a/regfile/regfile$10$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b329|t/a/regfile/reg0_b342  (
    .a({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_13 }),
    .b({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/ID_rs1$1$_placeOpt_13 }),
    .c({\t/a/ID_rs1$2$_placeOpt_4 ,\t/a/ID_rs1$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [9],\t/a/regfile/regfile$10$ [22]}),
    .e({\t/a/regfile/regfile$11$ [9],\t/a/regfile/regfile$11$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u351_o,_al_u708_o}),
    .q({\t/a/regfile/regfile$10$ [9],\t/a/regfile/regfile$10$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000011111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b330|t/a/regfile/reg0_b341  (
    .a({\t/a/ID_rs1$0$_placeOpt_11 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .b({\t/a/ID_rs1$1$_placeOpt_11 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$10$ [10],\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$2$_placeOpt_5 ,\t/a/regfile/regfile$10$ [21]}),
    .e({\t/a/regfile/regfile$11$ [10],\t/a/regfile/regfile$11$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u971_o,_al_u719_o}),
    .q({\t/a/regfile/regfile$10$ [10],\t/a/regfile/regfile$10$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000011111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b331|t/a/regfile/reg0_b340  (
    .a({\t/a/ID_rs1$0$_placeOpt_17 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .b({\t/a/ID_rs1$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$10$ [11],\t/a/ID_rs1$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$2$_placeOpt_3 ,\t/a/regfile/regfile$10$ [20]}),
    .e({\t/a/regfile/regfile$11$ [11],\t/a/regfile/regfile$11$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u960_o,_al_u750_o}),
    .q({\t/a/regfile/regfile$10$ [11],\t/a/regfile/regfile$10$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b332|t/a/regfile/reg0_b339  (
    .a({\t/a/ID_rs1$0$_placeOpt_17 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .b({\t/a/ID_rs1$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/ID_rs1$2$_placeOpt_3 ,\t/a/ID_rs1$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [12],\t/a/regfile/regfile$10$ [19]}),
    .e({\t/a/regfile/regfile$11$ [12],\t/a/regfile/regfile$11$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u929_o,_al_u782_o}),
    .q({\t/a/regfile/regfile$10$ [12],\t/a/regfile/regfile$10$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000011111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b333|t/a/regfile/reg0_b338  (
    .a({\t/a/ID_rs1$0$_placeOpt_11 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .b({\t/a/ID_rs1$1$_placeOpt_11 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$10$ [13],\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$2$_placeOpt_5 ,\t/a/regfile/regfile$10$ [18]}),
    .e({\t/a/regfile/regfile$11$ [13],\t/a/regfile/regfile$11$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u918_o,_al_u813_o}),
    .q({\t/a/regfile/regfile$10$ [13],\t/a/regfile/regfile$10$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000011111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b334|t/a/regfile/reg0_b337  (
    .a({\t/a/ID_rs1$0$_placeOpt_11 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .b({\t/a/ID_rs1$1$_placeOpt_11 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$10$ [14],\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$2$_placeOpt_5 ,\t/a/regfile/regfile$10$ [17]}),
    .e({\t/a/regfile/regfile$11$ [14],\t/a/regfile/regfile$11$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u887_o,_al_u824_o}),
    .q({\t/a/regfile/regfile$10$ [14],\t/a/regfile/regfile$10$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000011111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b335|t/a/regfile/reg0_b336  (
    .a({\t/a/ID_rs1$0$_placeOpt_9 ,\t/a/ID_rs1$0$_placeOpt_9 }),
    .b({\t/a/ID_rs1$1$_placeOpt_9 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .c({\t/a/regfile/regfile$10$ [15],\t/a/ID_rs1$2$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$2$_placeOpt_8 ,\t/a/regfile/regfile$10$ [16]}),
    .e({\t/a/regfile/regfile$11$ [15],\t/a/regfile/regfile$11$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u866_o,_al_u855_o}),
    .q({\t/a/regfile/regfile$10$ [15],\t/a/regfile/regfile$10$ [16]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b33|t/a/regfile/reg0_b63  (
    .a({\t/a/ID_rs1$0$_placeOpt_20 ,\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/a/ID_rs1$1$_placeOpt_20 ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/regfile/regfile$1$ [1],\t/a/regfile/regfile$0$ [31]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$0$ [1],\t/a/regfile/regfile$1$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u756_o,_al_u1199_o}),
    .q({\t/a/regfile/regfile$1$ [1],\t/a/regfile/regfile$1$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b34|t/a/regfile/reg0_b62  (
    .a({\t/a/ID_rs1$0$_placeOpt_10 ,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/ID_rs1$1$_placeOpt_10 ,\t/a/ID_rs2$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$0$ [2],\t/a/regfile/regfile$0$ [30]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [2],\t/a/regfile/regfile$1$ [30]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u525_o,_al_u1230_o}),
    .q({\t/a/regfile/regfile$1$ [2],\t/a/regfile/regfile$1$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*~D*C*B*A)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b352|t/a/regfile/reg0_b383  (
    .a({_al_u254_o,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2$1$_placeOpt_11 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$10$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$11$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b352_sel_is_3_o ,_al_u1204_o}),
    .q({\t/a/regfile/regfile$11$ [0],\t/a/regfile/regfile$11$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b353|t/a/regfile/reg0_b382  (
    .a({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/ID_rs2$2$_placeOpt_7 ,\t/a/ID_rs2$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [1],\t/a/regfile/regfile$10$ [30]}),
    .e({\t/a/regfile/regfile$11$ [1],\t/a/regfile/regfile$11$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1477_o,_al_u1235_o}),
    .q({\t/a/regfile/regfile$11$ [1],\t/a/regfile/regfile$11$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~A*~(B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~A*~(B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0001010100010001),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0101010101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b354|t/a/regfile/reg0_b381  (
    .a({\t/a/ID_rs2$2$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_11 }),
    .b({\t/a/ID_rs2$1$_placeOpt_9 ,\t/a/ID_rs2$1$_placeOpt_9 }),
    .c({\t/a/ID_rs2$0$_placeOpt_11 ,\t/a/ID_rs2$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [2],\t/a/regfile/regfile$10$ [29]}),
    .e({\t/a/regfile/regfile$11$ [2],\t/a/regfile/regfile$11$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1246_o,_al_u1267_o}),
    .q({\t/a/regfile/regfile$11$ [2],\t/a/regfile/regfile$11$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(A*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(A*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000101),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b355|t/a/regfile/reg0_b380  (
    .a({\t/a/ID_rs2$1$_placeOpt_20 ,\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2$1$_placeOpt_20 }),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [3],\t/a/regfile/regfile$10$ [28]}),
    .e({\t/a/regfile/regfile$11$ [3],\t/a/regfile/regfile$11$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1193_o,_al_u1298_o}),
    .q({\t/a/regfile/regfile$11$ [3],\t/a/regfile/regfile$11$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~B*~(C*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~B*~(C*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0001001100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0011001100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b356|t/a/regfile/reg0_b379  (
    .a({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/ID_rs2$2$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_12 }),
    .c({\t/a/ID_rs2$1$_placeOpt_12 ,\t/a/ID_rs2$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [4],\t/a/regfile/regfile$10$ [27]}),
    .e({\t/a/regfile/regfile$11$ [4],\t/a/regfile/regfile$11$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1162_o,_al_u1309_o}),
    .q({\t/a/regfile/regfile$11$ [4],\t/a/regfile/regfile$11$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~A*~(B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~A*~(B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0001010100010001),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0101010101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b357|t/a/regfile/reg0_b378  (
    .a({\t/a/ID_rs2$2$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_11 }),
    .b({\t/a/ID_rs2$1$_placeOpt_9 ,\t/a/ID_rs2$1$_placeOpt_9 }),
    .c({\t/a/ID_rs2$0$_placeOpt_11 ,\t/a/ID_rs2$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [5],\t/a/regfile/regfile$10$ [26]}),
    .e({\t/a/regfile/regfile$11$ [5],\t/a/regfile/regfile$11$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1141_o,_al_u1340_o}),
    .q({\t/a/regfile/regfile$11$ [5],\t/a/regfile/regfile$11$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b358|t/a/regfile/reg0_b377  (
    .a({\t/a/ID_rs2$0$_placeOpt_17 ,\t/a/ID_rs2$0$_placeOpt_17 }),
    .b({\t/a/ID_rs2$1$_placeOpt_8 ,\t/a/ID_rs2$1$_placeOpt_8 }),
    .c({\t/a/ID_rs2$2$_placeOpt_3 ,\t/a/ID_rs2$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [6],\t/a/regfile/regfile$10$ [25]}),
    .e({\t/a/regfile/regfile$11$ [6],\t/a/regfile/regfile$11$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1120_o,_al_u1351_o}),
    .q({\t/a/regfile/regfile$11$ [6],\t/a/regfile/regfile$11$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000011111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b359|t/a/regfile/reg0_b376  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2$1$_placeOpt_20 ,\t/a/ID_rs2$1$_placeOpt_20 }),
    .c({\t/a/regfile/regfile$10$ [7],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [2],\t/a/regfile/regfile$10$ [24]}),
    .e({\t/a/regfile/regfile$11$ [7],\t/a/regfile/regfile$11$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1099_o,_al_u1372_o}),
    .q({\t/a/regfile/regfile$11$ [7],\t/a/regfile/regfile$11$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b35|t/a/regfile/reg0_b61  (
    .a({\t/a/ID_rs2$0$_placeOpt_19 ,\t/a/ID_rs2$0$_placeOpt_19 }),
    .b({\t/a/ID_rs2$1$_placeOpt_19 ,\t/a/ID_rs2$1$_placeOpt_19 }),
    .c({\t/a/regfile/regfile$0$ [3],\t/a/regfile/regfile$0$ [29]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [3],\t/a/regfile/regfile$1$ [29]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1188_o,_al_u1262_o}),
    .q({\t/a/regfile/regfile$1$ [3],\t/a/regfile/regfile$1$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~A*~(B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~A*~(B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0001010100010001),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0101010101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b360|t/a/regfile/reg0_b375  (
    .a({\t/a/ID_rs2$2$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_11 }),
    .b({\t/a/ID_rs2$1$_placeOpt_9 ,\t/a/ID_rs2$1$_placeOpt_9 }),
    .c({\t/a/ID_rs2$0$_placeOpt_11 ,\t/a/ID_rs2$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [8],\t/a/regfile/regfile$10$ [23]}),
    .e({\t/a/regfile/regfile$11$ [8],\t/a/regfile/regfile$11$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1088_o,_al_u1403_o}),
    .q({\t/a/regfile/regfile$11$ [8],\t/a/regfile/regfile$11$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~B*~(C*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~B*~(C*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0001001100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0011001100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b361|t/a/regfile/reg0_b374  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2$2$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_12 }),
    .c({\t/a/ID_rs2$1$_placeOpt_12 ,\t/a/ID_rs2$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [9],\t/a/regfile/regfile$10$ [22]}),
    .e({\t/a/regfile/regfile$11$ [9],\t/a/regfile/regfile$11$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1057_o,_al_u1414_o}),
    .q({\t/a/regfile/regfile$11$ [9],\t/a/regfile/regfile$11$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b362|t/a/regfile/reg0_b373  (
    .a({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs2$0$_placeOpt_12 }),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_5 }),
    .c({\t/a/ID_rs2$2$_placeOpt_2 ,\t/a/ID_rs2$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [10],\t/a/regfile/regfile$10$ [21]}),
    .e({\t/a/regfile/regfile$11$ [10],\t/a/regfile/regfile$11$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1697_o,_al_u1445_o}),
    .q({\t/a/regfile/regfile$11$ [10],\t/a/regfile/regfile$11$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b363|t/a/regfile/reg0_b372  (
    .a({\t/a/ID_rs2$0$_placeOpt_13 ,\t/a/ID_rs2$0$_placeOpt_13 }),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs2$1$_placeOpt_17 }),
    .c({\t/a/ID_rs2$2$_placeOpt_3 ,\t/a/ID_rs2$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [11],\t/a/regfile/regfile$10$ [20]}),
    .e({\t/a/regfile/regfile$11$ [11],\t/a/regfile/regfile$11$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1666_o,_al_u1456_o}),
    .q({\t/a/regfile/regfile$11$ [11],\t/a/regfile/regfile$11$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000011111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b364|t/a/regfile/reg0_b371  (
    .a({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs2$0$_placeOpt_20 }),
    .b({\t/a/ID_rs2$1$_placeOpt_10 ,\t/a/ID_rs2$1$_placeOpt_10 }),
    .c({\t/a/regfile/regfile$10$ [12],\t/a/ID_rs2$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$2$_placeOpt_3 ,\t/a/regfile/regfile$10$ [19]}),
    .e({\t/a/regfile/regfile$11$ [12],\t/a/regfile/regfile$11$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1655_o,_al_u1498_o}),
    .q({\t/a/regfile/regfile$11$ [12],\t/a/regfile/regfile$11$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(A*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(A*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000101),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b365|t/a/regfile/reg0_b370  (
    .a({\t/a/ID_rs2$1$_placeOpt_8 ,\t/a/ID_rs2$0$_placeOpt_17 }),
    .b({\t/a/ID_rs2$0$_placeOpt_17 ,\t/a/ID_rs2$1$_placeOpt_8 }),
    .c({\t/a/ID_rs2$2$_placeOpt_2 ,\t/a/ID_rs2$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [13],\t/a/regfile/regfile$10$ [18]}),
    .e({\t/a/regfile/regfile$11$ [13],\t/a/regfile/regfile$11$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1624_o,_al_u1519_o}),
    .q({\t/a/regfile/regfile$11$ [13],\t/a/regfile/regfile$11$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(A*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(A*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000101),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b366|t/a/regfile/reg0_b369  (
    .a({\t/a/ID_rs2$1$_placeOpt_8 ,\t/a/ID_rs2$0$_placeOpt_17 }),
    .b({\t/a/ID_rs2$0$_placeOpt_17 ,\t/a/ID_rs2$1$_placeOpt_8 }),
    .c({\t/a/ID_rs2$2$_placeOpt_2 ,\t/a/ID_rs2$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [14],\t/a/regfile/regfile$10$ [17]}),
    .e({\t/a/regfile/regfile$11$ [14],\t/a/regfile/regfile$11$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1603_o,_al_u1550_o}),
    .q({\t/a/regfile/regfile$11$ [14],\t/a/regfile/regfile$11$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~A*~(B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~A*~(B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0001010100010001),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0101010101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b367|t/a/regfile/reg0_b368  (
    .a({\t/a/ID_rs2$2$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_20 }),
    .b({\t/a/ID_rs2$1$_placeOpt_10 ,\t/a/ID_rs2$1$_placeOpt_10 }),
    .c({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs2$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [15],\t/a/regfile/regfile$10$ [16]}),
    .e({\t/a/regfile/regfile$11$ [15],\t/a/regfile/regfile$11$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1592_o,_al_u1561_o}),
    .q({\t/a/regfile/regfile$11$ [15],\t/a/regfile/regfile$11$ [16]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b36|t/a/regfile/reg0_b60  (
    .a({\t/a/ID_rs1$0$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_16 }),
    .b({\t/a/ID_rs1$1$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$0$ [4],\t/a/regfile/regfile$0$ [28]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [4],\t/a/regfile/regfile$1$ [28]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u451_o,_al_u1293_o}),
    .q({\t/a/regfile/regfile$1$ [4],\t/a/regfile/regfile$1$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b37|t/a/regfile/reg0_b59  (
    .a({\t/a/ID_rs1$0$_placeOpt_10 ,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/ID_rs1$1$_placeOpt_10 ,\t/a/ID_rs2$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$0$ [5],\t/a/regfile/regfile$0$ [27]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [5],\t/a/regfile/regfile$1$ [27]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u420_o,_al_u1304_o}),
    .q({\t/a/regfile/regfile$1$ [5],\t/a/regfile/regfile$1$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b38|t/a/regfile/reg0_b58  (
    .a({\t/a/ID_rs1$0$_placeOpt_18 ,\t/a/ID_rs2$0$_placeOpt_20 }),
    .b({\t/a/ID_rs1$1$_placeOpt_18 ,\t/a/ID_rs2$1$_placeOpt_21 }),
    .c({\t/a/regfile/regfile$0$ [6],\t/a/regfile/regfile$0$ [26]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [6],\t/a/regfile/regfile$1$ [26]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u399_o,_al_u1335_o}),
    .q({\t/a/regfile/regfile$1$ [6],\t/a/regfile/regfile$1$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b39|t/a/regfile/reg0_b57  (
    .a({\t/a/ID_rs1$0$_placeOpt_14 ,\t/a/ID_rs2$0$_placeOpt_14 }),
    .b({\t/a/ID_rs1$1$_placeOpt_14 ,\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$1$ [7],\t/a/regfile/regfile$0$ [25]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$0$ [7],\t/a/regfile/regfile$1$ [25]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u388_o,_al_u1346_o}),
    .q({\t/a/regfile/regfile$1$ [7],\t/a/regfile/regfile$1$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b40|t/a/regfile/reg0_b56  (
    .a({\t/a/ID_rs1$0$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_16 }),
    .b({\t/a/ID_rs1$1$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_16 }),
    .c({\t/a/regfile/regfile$0$ [8],\t/a/regfile/regfile$0$ [24]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [8],\t/a/regfile/regfile$1$ [24]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u357_o,_al_u1367_o}),
    .q({\t/a/regfile/regfile$1$ [8],\t/a/regfile/regfile$1$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b41|t/a/regfile/reg0_b55  (
    .a({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/regfile/regfile$1$ [9],\t/a/regfile/regfile$0$ [23]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$0$ [9],\t/a/regfile/regfile$1$ [23]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u346_o,_al_u1398_o}),
    .q({\t/a/regfile/regfile$1$ [9],\t/a/regfile/regfile$1$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000000110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b42|t/a/regfile/reg0_b54  (
    .a({\t/a/regfile/regfile$0$ [10],\t/a/ID_rs2$0$_placeOpt_1 }),
    .b({\t/a/regfile/regfile$1$ [10],\t/a/ID_rs2$1$_placeOpt_16 }),
    .c({\t/a/ID_rs1$0$_placeOpt_3 ,\t/a/regfile/regfile$0$ [22]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_3 ,\t/a/regfile/regfile$1$ [22]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u966_o,_al_u1409_o}),
    .q({\t/a/regfile/regfile$1$ [10],\t/a/regfile/regfile$1$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000000110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b43|t/a/regfile/reg0_b53  (
    .a({\t/a/regfile/regfile$0$ [11],\t/a/ID_rs2$0$_placeOpt_12 }),
    .b({\t/a/regfile/regfile$1$ [11],\t/a/ID_rs2$1$_placeOpt_5 }),
    .c({\t/a/ID_rs1$0$_placeOpt_14 ,\t/a/regfile/regfile$0$ [21]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_14 ,\t/a/regfile/regfile$1$ [21]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u955_o,_al_u1440_o}),
    .q({\t/a/regfile/regfile$1$ [11],\t/a/regfile/regfile$1$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*D*C*~A*B)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*D*C*~A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b448|t/a/regfile/reg0_b479  (
    .a({\t/a/WB_rd [0],\t/a/ID_rs1$0$_placeOpt_16 }),
    .b({_al_u254_o,\t/a/ID_rs1$1$_placeOpt_16 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1$2$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$14$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$15$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b448_sel_is_3_o ,_al_u496_o}),
    .q({\t/a/regfile/regfile$14$ [0],\t/a/regfile/regfile$14$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111001100000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111101100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b449|t/a/regfile/reg0_b478  (
    .a({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/ID_rs1$0$_placeOpt_16 }),
    .b({\t/a/ID_rs1$1$_placeOpt_16 ,\t/a/ID_rs1$1$_placeOpt_16 }),
    .c({\t/a/regfile/regfile$14$ [1],\t/a/ID_rs1$2$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$2$_placeOpt_6 ,\t/a/regfile/regfile$14$ [30]}),
    .e({\t/a/regfile/regfile$15$ [1],\t/a/regfile/regfile$15$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u759_o,_al_u507_o}),
    .q({\t/a/regfile/regfile$14$ [1],\t/a/regfile/regfile$14$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000000110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b44|t/a/regfile/reg0_b52  (
    .a({\t/a/regfile/regfile$0$ [12],\t/a/ID_rs2$0$_placeOpt_20 }),
    .b({\t/a/regfile/regfile$1$ [12],\t/a/ID_rs2$1$_placeOpt_10 }),
    .c({\t/a/ID_rs1$0$_placeOpt_9 ,\t/a/regfile/regfile$0$ [20]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_9 ,\t/a/regfile/regfile$1$ [20]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u924_o,_al_u1451_o}),
    .q({\t/a/regfile/regfile$1$ [12],\t/a/regfile/regfile$1$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111001100000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111101100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b450|t/a/regfile/reg0_b477  (
    .a({\t/a/ID_rs1$0$_placeOpt_12 ,\t/a/ID_rs1$0$_placeOpt_12 }),
    .b({\t/a/ID_rs1$1$_placeOpt_12 ,\t/a/ID_rs1$1$_placeOpt_12 }),
    .c({\t/a/regfile/regfile$14$ [2],\t/a/ID_rs1$2$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$2$_placeOpt_8 ,\t/a/regfile/regfile$14$ [29]}),
    .e({\t/a/regfile/regfile$15$ [2],\t/a/regfile/regfile$15$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u528_o,_al_u559_o}),
    .q({\t/a/regfile/regfile$14$ [2],\t/a/regfile/regfile$14$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b451|t/a/regfile/reg0_b476  (
    .a({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_13 }),
    .b({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/ID_rs1$1$_placeOpt_13 }),
    .c({\t/a/ID_rs1$2$_placeOpt_4 ,\t/a/ID_rs1$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [3],\t/a/regfile/regfile$14$ [28]}),
    .e({\t/a/regfile/regfile$15$ [3],\t/a/regfile/regfile$15$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u465_o,_al_u570_o}),
    .q({\t/a/regfile/regfile$14$ [3],\t/a/regfile/regfile$14$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b452|t/a/regfile/reg0_b475  (
    .a({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_13 }),
    .b({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/ID_rs1$1$_placeOpt_13 }),
    .c({\t/a/ID_rs1$2$_placeOpt_4 ,\t/a/ID_rs1$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [4],\t/a/regfile/regfile$14$ [27]}),
    .e({\t/a/regfile/regfile$15$ [4],\t/a/regfile/regfile$15$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u454_o,_al_u601_o}),
    .q({\t/a/regfile/regfile$14$ [4],\t/a/regfile/regfile$14$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b453|t/a/regfile/reg0_b474  (
    .a({\t/a/ID_rs1$0$_placeOpt_9 ,\t/a/ID_rs1$0$_placeOpt_9 }),
    .b({\t/a/ID_rs1$1$_placeOpt_9 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .c({\t/a/ID_rs1$2$_placeOpt_3 ,\t/a/ID_rs1$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [5],\t/a/regfile/regfile$14$ [26]}),
    .e({\t/a/regfile/regfile$15$ [5],\t/a/regfile/regfile$15$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u423_o,_al_u612_o}),
    .q({\t/a/regfile/regfile$14$ [5],\t/a/regfile/regfile$14$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111001100000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111101100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b454|t/a/regfile/reg0_b473  (
    .a({\t/a/ID_rs1$0$_placeOpt_17 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .b({\t/a/ID_rs1$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$14$ [6],\t/a/ID_rs1$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$2$_placeOpt_3 ,\t/a/regfile/regfile$14$ [25]}),
    .e({\t/a/regfile/regfile$15$ [6],\t/a/regfile/regfile$15$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u402_o,_al_u633_o}),
    .q({\t/a/regfile/regfile$14$ [6],\t/a/regfile/regfile$14$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(B*~(D*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(B*~(D*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0100000011001100),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1100100011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b455|t/a/regfile/reg0_b472  (
    .a({\t/a/ID_rs1$0$_placeOpt_1 ,\t/a/ID_rs1$0$_placeOpt_1 }),
    .b({\t/a/ID_rs1$2$_placeOpt_1 ,\t/a/ID_rs1$1$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$14$ [7],\t/a/ID_rs1$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_1 ,\t/a/regfile/regfile$14$ [24]}),
    .e({\t/a/regfile/regfile$15$ [7],\t/a/regfile/regfile$15$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u391_o,_al_u654_o}),
    .q({\t/a/regfile/regfile$14$ [7],\t/a/regfile/regfile$14$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b456|t/a/regfile/reg0_b471  (
    .a({\t/a/ID_rs1$0$_placeOpt_12 ,\t/a/ID_rs1$0$_placeOpt_12 }),
    .b({\t/a/ID_rs1$1$_placeOpt_12 ,\t/a/ID_rs1$1$_placeOpt_12 }),
    .c({\t/a/ID_rs1$2$_placeOpt_8 ,\t/a/ID_rs1$2$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [8],\t/a/regfile/regfile$14$ [23]}),
    .e({\t/a/regfile/regfile$15$ [8],\t/a/regfile/regfile$15$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u360_o,_al_u675_o}),
    .q({\t/a/regfile/regfile$14$ [8],\t/a/regfile/regfile$14$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111001100000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111101100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b457|t/a/regfile/reg0_b470  (
    .a({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_13 }),
    .b({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/ID_rs1$1$_placeOpt_13 }),
    .c({\t/a/regfile/regfile$14$ [9],\t/a/ID_rs1$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$2$_placeOpt_4 ,\t/a/regfile/regfile$14$ [22]}),
    .e({\t/a/regfile/regfile$15$ [9],\t/a/regfile/regfile$15$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u349_o,_al_u706_o}),
    .q({\t/a/regfile/regfile$14$ [9],\t/a/regfile/regfile$14$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b458|t/a/regfile/reg0_b469  (
    .a({\t/a/ID_rs1$0$_placeOpt_11 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .b({\t/a/ID_rs1$1$_placeOpt_11 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/ID_rs1$2$_placeOpt_5 ,\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [10],\t/a/regfile/regfile$14$ [21]}),
    .e({\t/a/regfile/regfile$15$ [10],\t/a/regfile/regfile$15$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u969_o,_al_u717_o}),
    .q({\t/a/regfile/regfile$14$ [10],\t/a/regfile/regfile$14$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b459|t/a/regfile/reg0_b468  (
    .a({\t/a/ID_rs1$0$_placeOpt_21 ,\t/a/ID_rs1$0$_placeOpt_21 }),
    .b({\t/a/ID_rs1$1$_placeOpt_21 ,\t/a/ID_rs1$1$_placeOpt_21 }),
    .c({\t/a/ID_rs1$2$_placeOpt_3 ,\t/a/ID_rs1$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [11],\t/a/regfile/regfile$14$ [20]}),
    .e({\t/a/regfile/regfile$15$ [11],\t/a/regfile/regfile$15$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u958_o,_al_u748_o}),
    .q({\t/a/regfile/regfile$14$ [11],\t/a/regfile/regfile$14$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000000110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b45|t/a/regfile/reg0_b51  (
    .a({\t/a/regfile/regfile$0$ [13],\t/a/ID_rs2$0$_placeOpt_18 }),
    .b({\t/a/regfile/regfile$1$ [13],\t/a/ID_rs2$1$_placeOpt_19 }),
    .c({\t/a/ID_rs1$0$_placeOpt_14 ,\t/a/regfile/regfile$0$ [19]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_14 ,\t/a/regfile/regfile$1$ [19]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u913_o,_al_u1493_o}),
    .q({\t/a/regfile/regfile$1$ [13],\t/a/regfile/regfile$1$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b460|t/a/regfile/reg0_b467  (
    .a({\t/a/ID_rs1$0$_placeOpt_17 ,\t/a/ID_rs1$0$_placeOpt_17 }),
    .b({\t/a/ID_rs1$1$_placeOpt_17 ,\t/a/ID_rs1$1$_placeOpt_17 }),
    .c({\t/a/ID_rs1$2$_placeOpt_3 ,\t/a/ID_rs1$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [12],\t/a/regfile/regfile$14$ [19]}),
    .e({\t/a/regfile/regfile$15$ [12],\t/a/regfile/regfile$15$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u927_o,_al_u780_o}),
    .q({\t/a/regfile/regfile$14$ [12],\t/a/regfile/regfile$14$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b461|t/a/regfile/reg0_b466  (
    .a({\t/a/ID_rs1$0$_placeOpt_21 ,\t/a/ID_rs1$0$_placeOpt_21 }),
    .b({\t/a/ID_rs1$1$_placeOpt_21 ,\t/a/ID_rs1$1$_placeOpt_21 }),
    .c({\t/a/ID_rs1$2$_placeOpt_3 ,\t/a/ID_rs1$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [13],\t/a/regfile/regfile$14$ [18]}),
    .e({\t/a/regfile/regfile$15$ [13],\t/a/regfile/regfile$15$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u916_o,_al_u811_o}),
    .q({\t/a/regfile/regfile$14$ [13],\t/a/regfile/regfile$14$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111001100000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111101100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b462|t/a/regfile/reg0_b465  (
    .a({\t/a/ID_rs1$0$_placeOpt_11 ,\t/a/ID_rs1$0$_placeOpt_11 }),
    .b({\t/a/ID_rs1$1$_placeOpt_11 ,\t/a/ID_rs1$1$_placeOpt_11 }),
    .c({\t/a/regfile/regfile$14$ [14],\t/a/ID_rs1$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$2$_placeOpt_5 ,\t/a/regfile/regfile$14$ [17]}),
    .e({\t/a/regfile/regfile$15$ [14],\t/a/regfile/regfile$15$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u885_o,_al_u822_o}),
    .q({\t/a/regfile/regfile$14$ [14],\t/a/regfile/regfile$14$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b463|t/a/regfile/reg0_b464  (
    .a({\t/a/ID_rs1$0$_placeOpt_9 ,\t/a/ID_rs1$0$_placeOpt_9 }),
    .b({\t/a/ID_rs1$1$_placeOpt_9 ,\t/a/ID_rs1$1$_placeOpt_9 }),
    .c({\t/a/ID_rs1$2$_placeOpt_3 ,\t/a/ID_rs1$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [15],\t/a/regfile/regfile$14$ [16]}),
    .e({\t/a/regfile/regfile$15$ [15],\t/a/regfile/regfile$15$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u864_o,_al_u853_o}),
    .q({\t/a/regfile/regfile$14$ [15],\t/a/regfile/regfile$14$ [16]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000000110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b46|t/a/regfile/reg0_b50  (
    .a({\t/a/regfile/regfile$0$ [14],\t/a/ID_rs2$0$_placeOpt_9 }),
    .b({\t/a/regfile/regfile$1$ [14],\t/a/ID_rs2$1$_placeOpt_17 }),
    .c({\t/a/ID_rs1$0$_placeOpt_21 ,\t/a/regfile/regfile$0$ [18]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_21 ,\t/a/regfile/regfile$1$ [18]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u882_o,_al_u1514_o}),
    .q({\t/a/regfile/regfile$1$ [14],\t/a/regfile/regfile$1$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*D*C*A*B)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*D*C*A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b480|t/a/regfile/reg0_b511  (
    .a({\t/a/WB_rd [0],\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({_al_u254_o,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$14$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$15$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b480_sel_is_3_o ,_al_u1202_o}),
    .q({\t/a/regfile/regfile$15$ [0],\t/a/regfile/regfile$15$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b481|t/a/regfile/reg0_b510  (
    .a({\t/a/ID_rs2$0$_placeOpt_21 ,\t/a/ID_rs2$0$_placeOpt_21 }),
    .b({\t/a/ID_rs2$1$_placeOpt_15 ,\t/a/ID_rs2$1$_placeOpt_15 }),
    .c({\t/a/ID_rs2$2$_placeOpt_7 ,\t/a/ID_rs2$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [1],\t/a/regfile/regfile$14$ [30]}),
    .e({\t/a/regfile/regfile$15$ [1],\t/a/regfile/regfile$15$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1475_o,_al_u1233_o}),
    .q({\t/a/regfile/regfile$15$ [1],\t/a/regfile/regfile$15$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(A*~(C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(A*~(C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0010101000001010),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1010101010001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b482|t/a/regfile/reg0_b509  (
    .a({\t/a/ID_rs2$2$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_15 }),
    .b({\t/a/ID_rs2$0$_placeOpt_15 ,\t/a/ID_rs2$1$_placeOpt_9 }),
    .c({\t/a/ID_rs2$1$_placeOpt_9 ,\t/a/ID_rs2$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [2],\t/a/regfile/regfile$14$ [29]}),
    .e({\t/a/regfile/regfile$15$ [2],\t/a/regfile/regfile$15$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1244_o,_al_u1265_o}),
    .q({\t/a/regfile/regfile$15$ [2],\t/a/regfile/regfile$15$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b483|t/a/regfile/reg0_b508  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2$2$_placeOpt_10 ,\t/a/ID_rs2$2$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [3],\t/a/regfile/regfile$14$ [28]}),
    .e({\t/a/regfile/regfile$15$ [3],\t/a/regfile/regfile$15$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1191_o,_al_u1296_o}),
    .q({\t/a/regfile/regfile$15$ [3],\t/a/regfile/regfile$15$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(A*~(B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(A*~(B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0010101000100010),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1010101010100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b484|t/a/regfile/reg0_b507  (
    .a({\t/a/ID_rs2$2$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/ID_rs2$1$_placeOpt_12 ,\t/a/ID_rs2$1$_placeOpt_12 }),
    .c({\t/a/ID_rs2$0$_placeOpt_22 ,\t/a/ID_rs2$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [4],\t/a/regfile/regfile$14$ [27]}),
    .e({\t/a/regfile/regfile$15$ [4],\t/a/regfile/regfile$15$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1160_o,_al_u1307_o}),
    .q({\t/a/regfile/regfile$15$ [4],\t/a/regfile/regfile$15$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(B*~(C*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(B*~(C*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0100110000001100),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1100110010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b485|t/a/regfile/reg0_b506  (
    .a({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs2$0$_placeOpt_20 }),
    .b({\t/a/ID_rs2$2$_placeOpt_4 ,\t/a/ID_rs2$1$_placeOpt_21 }),
    .c({\t/a/ID_rs2$1$_placeOpt_21 ,\t/a/ID_rs2$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [5],\t/a/regfile/regfile$14$ [26]}),
    .e({\t/a/regfile/regfile$15$ [5],\t/a/regfile/regfile$15$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1139_o,_al_u1338_o}),
    .q({\t/a/regfile/regfile$15$ [5],\t/a/regfile/regfile$15$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b486|t/a/regfile/reg0_b505  (
    .a({\t/a/ID_rs2$0$_placeOpt_9 ,\t/a/ID_rs2$0$_placeOpt_9 }),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs2$1$_placeOpt_17 }),
    .c({\t/a/ID_rs2$2$_placeOpt_3 ,\t/a/ID_rs2$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [6],\t/a/regfile/regfile$14$ [25]}),
    .e({\t/a/regfile/regfile$15$ [6],\t/a/regfile/regfile$15$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1118_o,_al_u1349_o}),
    .q({\t/a/regfile/regfile$15$ [6],\t/a/regfile/regfile$15$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b487|t/a/regfile/reg0_b504  (
    .a({\t/a/ID_rs2$0$_placeOpt_10 ,\t/a/ID_rs2$0$_placeOpt_10 }),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2$2$_placeOpt_10 ,\t/a/ID_rs2$2$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [7],\t/a/regfile/regfile$14$ [24]}),
    .e({\t/a/regfile/regfile$15$ [7],\t/a/regfile/regfile$15$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1097_o,_al_u1370_o}),
    .q({\t/a/regfile/regfile$15$ [7],\t/a/regfile/regfile$15$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(B*~(A*~(C*~(0)*~(D)+C*0*~(D)+~(C)*0*D+C*0*D)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(B*~(A*~(C*~(1)*~(D)+C*1*~(D)+~(C)*1*D+C*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0100010011000100),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1100110011000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b488|t/a/regfile/reg0_b503  (
    .a({\t/a/ID_rs2$1$_placeOpt_9 ,\t/a/ID_rs2$0$_placeOpt_11 }),
    .b({\t/a/ID_rs2$2$_placeOpt_4 ,\t/a/ID_rs2$1$_placeOpt_9 }),
    .c({\t/a/regfile/regfile$14$ [8],\t/a/ID_rs2$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_11 ,\t/a/regfile/regfile$14$ [23]}),
    .e({\t/a/regfile/regfile$15$ [8],\t/a/regfile/regfile$15$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1086_o,_al_u1401_o}),
    .q({\t/a/regfile/regfile$15$ [8],\t/a/regfile/regfile$15$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(A*~(B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(A*~(B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0010101000100010),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1010101010100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b489|t/a/regfile/reg0_b502  (
    .a({\t/a/ID_rs2$2$_placeOpt_5 ,\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2$1$_placeOpt_12 ,\t/a/ID_rs2$1$_placeOpt_12 }),
    .c({\t/a/ID_rs2 [0],\t/a/ID_rs2$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [9],\t/a/regfile/regfile$14$ [22]}),
    .e({\t/a/regfile/regfile$15$ [9],\t/a/regfile/regfile$15$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1055_o,_al_u1412_o}),
    .q({\t/a/regfile/regfile$15$ [9],\t/a/regfile/regfile$15$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b490|t/a/regfile/reg0_b501  (
    .a({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs2$0$_placeOpt_12 }),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_5 }),
    .c({\t/a/ID_rs2$2$_placeOpt_2 ,\t/a/ID_rs2$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [10],\t/a/regfile/regfile$14$ [21]}),
    .e({\t/a/regfile/regfile$15$ [10],\t/a/regfile/regfile$15$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1695_o,_al_u1443_o}),
    .q({\t/a/regfile/regfile$15$ [10],\t/a/regfile/regfile$15$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111001100000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111101100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b491|t/a/regfile/reg0_b500  (
    .a({\t/a/ID_rs2$0$_placeOpt_9 ,\t/a/ID_rs2$0$_placeOpt_9 }),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs2$1$_placeOpt_17 }),
    .c({\t/a/regfile/regfile$14$ [11],\t/a/ID_rs2$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$2$_placeOpt_3 ,\t/a/regfile/regfile$14$ [20]}),
    .e({\t/a/regfile/regfile$15$ [11],\t/a/regfile/regfile$15$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1664_o,_al_u1454_o}),
    .q({\t/a/regfile/regfile$15$ [11],\t/a/regfile/regfile$15$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b492|t/a/regfile/reg0_b499  (
    .a({\t/a/ID_rs2$0$_placeOpt_13 ,\t/a/ID_rs2$0$_placeOpt_13 }),
    .b({\t/a/ID_rs2$1$_placeOpt_17 ,\t/a/ID_rs2$1$_placeOpt_17 }),
    .c({\t/a/ID_rs2$2$_placeOpt_3 ,\t/a/ID_rs2$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [12],\t/a/regfile/regfile$14$ [19]}),
    .e({\t/a/regfile/regfile$15$ [12],\t/a/regfile/regfile$15$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1653_o,_al_u1496_o}),
    .q({\t/a/regfile/regfile$15$ [12],\t/a/regfile/regfile$15$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b493|t/a/regfile/reg0_b498  (
    .a({\t/a/ID_rs2$0$_placeOpt_9 ,\t/a/ID_rs2$0$_placeOpt_9 }),
    .b({\t/a/ID_rs2$1$_placeOpt_14 ,\t/a/ID_rs2$1$_placeOpt_14 }),
    .c({\t/a/ID_rs2$2$_placeOpt_3 ,\t/a/ID_rs2$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [13],\t/a/regfile/regfile$14$ [18]}),
    .e({\t/a/regfile/regfile$15$ [13],\t/a/regfile/regfile$15$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1622_o,_al_u1517_o}),
    .q({\t/a/regfile/regfile$15$ [13],\t/a/regfile/regfile$15$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(A*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(A*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000001010000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b494|t/a/regfile/reg0_b497  (
    .a({\t/a/ID_rs2$1$_placeOpt_8 ,\t/a/ID_rs2$0$_placeOpt_17 }),
    .b({\t/a/ID_rs2$0$_placeOpt_17 ,\t/a/ID_rs2$1$_placeOpt_8 }),
    .c({\t/a/ID_rs2$2$_placeOpt_2 ,\t/a/ID_rs2$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [14],\t/a/regfile/regfile$14$ [17]}),
    .e({\t/a/regfile/regfile$15$ [14],\t/a/regfile/regfile$15$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1601_o,_al_u1548_o}),
    .q({\t/a/regfile/regfile$15$ [14],\t/a/regfile/regfile$15$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111001100000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111101100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b495|t/a/regfile/reg0_b496  (
    .a({\t/a/ID_rs2$0$_placeOpt_20 ,\t/a/ID_rs2$0$_placeOpt_20 }),
    .b({\t/a/ID_rs2$1$_placeOpt_10 ,\t/a/ID_rs2$1$_placeOpt_10 }),
    .c({\t/a/regfile/regfile$14$ [15],\t/a/ID_rs2$2$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$2$_placeOpt_3 ,\t/a/regfile/regfile$14$ [16]}),
    .e({\t/a/regfile/regfile$15$ [15],\t/a/regfile/regfile$15$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1590_o,_al_u1559_o}),
    .q({\t/a/regfile/regfile$15$ [15],\t/a/regfile/regfile$15$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b512|t/a/regfile/reg0_b543  (
    .a({_al_u256_o,_al_u488_o}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1$0$_placeOpt_10 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1$1$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$16$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$17$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b512_sel_is_3_o ,_al_u489_o}),
    .q({\t/a/regfile/regfile$16$ [0],\t/a/regfile/regfile$16$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*~B*~D*C+~A*~B*D*C"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("A*~B*~D*~C+A*~B*D*~C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0001001100010011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b513|t/a/regfile/reg0_b541  (
    .a({\t/a/ID_rs1$0$_placeOpt_5 ,_al_u551_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_5 ,\t/a/ID_rs1$0$_placeOpt_5 }),
    .c({\t/a/regfile/regfile$17$ [1],\t/a/ID_rs1$1$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({open_n37987,\t/a/regfile/regfile$16$ [29]}),
    .e({\t/a/regfile/regfile$16$ [1],\t/a/regfile/regfile$17$ [29]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u766_o,_al_u552_o}),
    .q({\t/a/regfile/regfile$16$ [1],\t/a/regfile/regfile$16$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~A*~D*~B*~C+~A*D*~B*~C+~A*~D*B*~C+~A*D*B*~C+~A*~D*~B*C+~A*~D*B*C"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~A*D*~B*~C+~A*D*B*~C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000010101010101),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b514|t/a/regfile/reg0_b539  (
    .a({\t/a/ID_rs1$1$_placeOpt_7 ,_al_u593_o}),
    .b({open_n38003,\t/a/ID_rs1$0$_placeOpt_7 }),
    .c({\t/a/regfile/regfile$17$ [2],\t/a/ID_rs1$1$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_7 ,\t/a/regfile/regfile$16$ [27]}),
    .e({\t/a/regfile/regfile$16$ [2],\t/a/regfile/regfile$17$ [27]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u535_o,_al_u594_o}),
    .q({\t/a/regfile/regfile$16$ [2],\t/a/regfile/regfile$16$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~C*~A*~D*~B+C*~A*~D*~B+C*~A*D*~B+~C*~A*~D*B+C*~A*~D*B+C*~A*D*B"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~C*~A*~D*~B+~C*~A*~D*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0101000001010101),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b515|t/a/regfile/reg0_b534  (
    .a({\t/a/ID_rs1$1$_placeOpt_8 ,_al_u698_o}),
    .b({open_n38019,\t/a/ID_rs1$0$_placeOpt_8 }),
    .c({\t/a/ID_rs1$0$_placeOpt_8 ,\t/a/ID_rs1$1$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$16$ [3],\t/a/regfile/regfile$16$ [22]}),
    .e({\t/a/regfile/regfile$17$ [3],\t/a/regfile/regfile$17$ [22]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u472_o,_al_u699_o}),
    .q({\t/a/regfile/regfile$16$ [3],\t/a/regfile/regfile$16$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b516|t/a/regfile/reg0_b532  (
    .a({_al_u446_o,_al_u740_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$16$ [4],\t/a/regfile/regfile$16$ [20]}),
    .e({\t/a/regfile/regfile$17$ [4],\t/a/regfile/regfile$17$ [20]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u447_o,_al_u741_o}),
    .q({\t/a/regfile/regfile$16$ [4],\t/a/regfile/regfile$16$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~C*~B*~A*~D+C*~B*~A*~D+~C*~B*A*~D+C*~B*A*~D+~C*~B*~A*D+~C*~B*A*D"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("C*~B*~A*~D+C*~B*A*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001100110011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b517|t/a/regfile/reg0_b530  (
    .a({open_n38050,_al_u803_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .c({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [5],\t/a/regfile/regfile$16$ [18]}),
    .e({\t/a/regfile/regfile$16$ [5],\t/a/regfile/regfile$17$ [18]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u430_o,_al_u804_o}),
    .q({\t/a/regfile/regfile$16$ [5],\t/a/regfile/regfile$16$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*~B*~C*D+~A*~B*C*D"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("A*~B*~C*~D+A*~B*C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0001000100110011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b518|t/a/regfile/reg0_b528  (
    .a({\t/a/ID_rs1$0$_placeOpt_14 ,_al_u845_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_14 ,\t/a/ID_rs1$0$_placeOpt_14 }),
    .c({open_n38066,\t/a/ID_rs1$1$_placeOpt_14 }),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [6],\t/a/regfile/regfile$16$ [16]}),
    .e({\t/a/regfile/regfile$16$ [6],\t/a/regfile/regfile$17$ [16]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u409_o,_al_u846_o}),
    .q({\t/a/regfile/regfile$16$ [6],\t/a/regfile/regfile$16$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(B*~(~A*~(C*~(0)*~(D)+C*0*~(D)+~(C)*0*D+C*0*D)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(B*~(~A*~(C*~(1)*~(D)+C*1*~(D)+~(C)*1*D+C*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1000100011001000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1100110011001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b519|t/a/regfile/reg0_b525  (
    .a({\t/a/ID_rs1$1$_placeOpt_7 ,_al_u908_o}),
    .b({_al_u383_o,\t/a/ID_rs1$0$_placeOpt_7 }),
    .c({\t/a/regfile/regfile$16$ [7],\t/a/ID_rs1$1$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_7 ,\t/a/regfile/regfile$16$ [13]}),
    .e({\t/a/regfile/regfile$17$ [7],\t/a/regfile/regfile$17$ [13]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u384_o,_al_u909_o}),
    .q({\t/a/regfile/regfile$16$ [7],\t/a/regfile/regfile$16$ [13]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~B*~C*~D*~A+B*~C*~D*~A+B*~C*D*~A+~B*~C*~D*A+B*~C*~D*A+B*~C*D*A"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~B*~C*~D*~A+~B*~C*~D*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000110000001111),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b520|t/a/regfile/reg0_b523  (
    .a({open_n38097,_al_u950_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .c({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/ID_rs1$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$16$ [8],\t/a/regfile/regfile$16$ [11]}),
    .e({\t/a/regfile/regfile$17$ [8],\t/a/regfile/regfile$17$ [11]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u367_o,_al_u951_o}),
    .q({\t/a/regfile/regfile$16$ [8],\t/a/regfile/regfile$16$ [11]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*~B*C*D"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b522|t/a/regfile/reg0_b521  (
    .a({\t/a/ID_rs1$0$_placeOpt_8 ,_al_u341_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_8 ,\t/a/ID_rs1$0$_placeOpt_8 }),
    .c({\t/a/regfile/regfile$16$ [10],\t/a/ID_rs1$1$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({open_n38113,\t/a/regfile/regfile$16$ [9]}),
    .e(\t/a/regfile/regfile$17$ [10:9]),
    .mi(\t/a/reg_writedat [10:9]),
    .sr(rst_pad),
    .f({_al_u976_o,_al_u342_o}),
    .q(\t/a/regfile/regfile$16$ [10:9]));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b524|t/a/regfile/reg0_b542  (
    .a({\t/a/ID_rs1$0$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_2 }),
    .b({\t/a/regfile/regfile$16$ [12],\t/a/ID_rs1$1$_placeOpt_2 }),
    .c({\t/a/ID_rs1$1$_placeOpt_2 ,\t/a/regfile/regfile$16$ [30]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [12],\t/a/regfile/regfile$17$ [30]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u934_o,_al_u514_o}),
    .q({\t/a/regfile/regfile$16$ [12],\t/a/regfile/regfile$16$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b526|t/a/regfile/reg0_b540  (
    .a({\t/a/ID_rs1$0$_placeOpt_8 ,\t/a/ID_rs1$0$_placeOpt_8 }),
    .b({\t/a/ID_rs1$1$_placeOpt_8 ,\t/a/ID_rs1$1$_placeOpt_8 }),
    .c({\t/a/regfile/regfile$16$ [14],\t/a/regfile/regfile$16$ [28]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [14],\t/a/regfile/regfile$17$ [28]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u892_o,_al_u577_o}),
    .q({\t/a/regfile/regfile$16$ [14],\t/a/regfile/regfile$16$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b527|t/a/regfile/reg0_b538  (
    .a({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/regfile/regfile$16$ [15],\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/regfile/regfile$16$ [26]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [15],\t/a/regfile/regfile$17$ [26]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u871_o,_al_u619_o}),
    .q({\t/a/regfile/regfile$16$ [15],\t/a/regfile/regfile$16$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b529|t/a/regfile/reg0_b537  (
    .a({\t/a/regfile/regfile$16$ [17],\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/regfile/regfile$16$ [25]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [17],\t/a/regfile/regfile$17$ [25]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u829_o,_al_u640_o}),
    .q({\t/a/regfile/regfile$16$ [17],\t/a/regfile/regfile$16$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b531|t/a/regfile/reg0_b536  (
    .a({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/regfile/regfile$17$ [19],\t/a/regfile/regfile$16$ [24]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$16$ [19],\t/a/regfile/regfile$17$ [24]}),
    .mi({\t/a/reg_writedat [19],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u787_o,_al_u661_o}),
    .q({\t/a/regfile/regfile$16$ [19],\t/a/regfile/regfile$16$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b533|t/a/regfile/reg0_b535  (
    .a({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/regfile/regfile$16$ [21],\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/regfile/regfile$16$ [23]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [21],\t/a/regfile/regfile$17$ [23]}),
    .mi({\t/a/reg_writedat [21],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u724_o,_al_u682_o}),
    .q({\t/a/regfile/regfile$16$ [21],\t/a/regfile/regfile$16$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*~D*~C*A*B)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*~D*~C*A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b544|t/a/regfile/reg0_b574  (
    .a({\t/a/WB_rd [0],_al_u1225_o}),
    .b({_al_u256_o,\t/a/ID_rs2$0$_placeOpt_22 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2$1$_placeOpt_11 }),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$16$ [30]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$17$ [30]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b544_sel_is_3_o ,_al_u1226_o}),
    .q({\t/a/regfile/regfile$17$ [0],\t/a/regfile/regfile$17$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*~D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*~D*C*B"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("A*~D*~C*~B+A*~D*~C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000001011111),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b545|t/a/regfile/reg0_b572  (
    .a({\t/a/ID_rs2$0$_placeOpt_4 ,_al_u1288_o}),
    .b({open_n38222,\t/a/ID_rs2$0$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$17$ [1],\t/a/ID_rs2$1$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_1 ,\t/a/regfile/regfile$16$ [28]}),
    .e({\t/a/regfile/regfile$16$ [1],\t/a/regfile/regfile$17$ [28]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1482_o,_al_u1289_o}),
    .q({\t/a/regfile/regfile$17$ [1],\t/a/regfile/regfile$17$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001100000011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b546|t/a/regfile/reg0_b570  (
    .a({open_n38238,_al_u1330_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$16$ [2],\t/a/ID_rs2$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [2],\t/a/regfile/regfile$16$ [26]}),
    .e({\t/a/ID_rs2$0$_placeOpt_2 ,\t/a/regfile/regfile$17$ [26]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1251_o,_al_u1331_o}),
    .q({\t/a/regfile/regfile$17$ [2],\t/a/regfile/regfile$17$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b547|t/a/regfile/reg0_b567  (
    .a({_al_u1183_o,_al_u1393_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_7 ,\t/a/ID_rs2$0$_placeOpt_7 }),
    .c({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/ID_rs2$1$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$16$ [3],\t/a/regfile/regfile$16$ [23]}),
    .e({\t/a/regfile/regfile$17$ [3],\t/a/regfile/regfile$17$ [23]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1184_o,_al_u1394_o}),
    .q({\t/a/regfile/regfile$17$ [3],\t/a/regfile/regfile$17$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+~A*B*~C*D"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000010110101111),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b548|t/a/regfile/reg0_b565  (
    .a({\t/a/ID_rs2$0$_placeOpt_7 ,_al_u1435_o}),
    .b({open_n38269,\t/a/ID_rs2$0$_placeOpt_7 }),
    .c({\t/a/regfile/regfile$16$ [4],\t/a/ID_rs2$1$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [4],\t/a/regfile/regfile$16$ [21]}),
    .e({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/regfile/regfile$17$ [21]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1167_o,_al_u1436_o}),
    .q({\t/a/regfile/regfile$17$ [4],\t/a/regfile/regfile$17$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+D*~B*C*A"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~D*~B*~C*~A+~D*~B*~C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b549|t/a/regfile/reg0_b561  (
    .a({open_n38285,_al_u1540_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_6 }),
    .c({\t/a/regfile/regfile$16$ [5],\t/a/ID_rs2$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_6 ,\t/a/regfile/regfile$16$ [17]}),
    .e({\t/a/regfile/regfile$17$ [5],\t/a/regfile/regfile$17$ [17]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1146_o,_al_u1541_o}),
    .q({\t/a/regfile/regfile$17$ [5],\t/a/regfile/regfile$17$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~A*~D*~B*~C+A*~D*~B*~C+~A*~D*B*~C+A*~D*B*~C+~A*~D*~B*C+~A*~D*B*C"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("A*~D*~B*~C+A*~D*B*~C"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000001011111),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b550|t/a/regfile/reg0_b559  (
    .a({\t/a/ID_rs2$0$_placeOpt_18 ,_al_u1582_o}),
    .b({open_n38301,\t/a/ID_rs2$0$_placeOpt_18 }),
    .c({\t/a/regfile/regfile$17$ [6],\t/a/ID_rs2$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/regfile/regfile$16$ [15]}),
    .e({\t/a/regfile/regfile$16$ [6],\t/a/regfile/regfile$17$ [15]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1125_o,_al_u1583_o}),
    .q({\t/a/regfile/regfile$17$ [6],\t/a/regfile/regfile$17$ [15]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~C*~B*~D*~A+C*~B*~D*~A+C*~B*D*~A+~C*~B*~D*A+C*~B*~D*A+C*~B*D*A"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~C*~B*~D*~A+~C*~B*~D*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b551|t/a/regfile/reg0_b556  (
    .a({open_n38317,_al_u1645_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .c({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$16$ [7],\t/a/regfile/regfile$16$ [12]}),
    .e({\t/a/regfile/regfile$17$ [7],\t/a/regfile/regfile$17$ [12]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1104_o,_al_u1646_o}),
    .q({\t/a/regfile/regfile$17$ [7],\t/a/regfile/regfile$17$ [12]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b552|t/a/regfile/reg0_b554  (
    .a({_al_u1078_o,_al_u1687_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$16$ [8],\t/a/ID_rs2$1$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/regfile/regfile$16$ [10]}),
    .e({\t/a/regfile/regfile$17$ [8],\t/a/regfile/regfile$17$ [10]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1079_o,_al_u1688_o}),
    .q({\t/a/regfile/regfile$17$ [8],\t/a/regfile/regfile$17$ [10]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b553|t/a/regfile/reg0_b575  (
    .a({\t/a/regfile/regfile$17$ [9],\t/a/ID_rs2$0$_placeOpt_4 }),
    .b({\t/a/regfile/regfile$16$ [9],\t/a/ID_rs2$1$_placeOpt_3 }),
    .c({\t/a/ID_rs2$1$_placeOpt_3 ,\t/a/regfile/regfile$16$ [31]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/regfile/regfile$17$ [31]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1062_o,_al_u1209_o}),
    .q({\t/a/regfile/regfile$17$ [9],\t/a/regfile/regfile$17$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b555|t/a/regfile/reg0_b573  (
    .a({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$16$ [11],\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/regfile/regfile$16$ [29]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [11],\t/a/regfile/regfile$17$ [29]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1671_o,_al_u1272_o}),
    .q({\t/a/regfile/regfile$17$ [11],\t/a/regfile/regfile$17$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001100010001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b557|t/a/regfile/reg0_b571  (
    .a({\t/a/regfile/regfile$16$ [13],\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/regfile/regfile$17$ [13],\t/a/regfile/regfile$16$ [27]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/regfile/regfile$17$ [27]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1629_o,_al_u1314_o}),
    .q({\t/a/regfile/regfile$17$ [13],\t/a/regfile/regfile$17$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b558|t/a/regfile/reg0_b569  (
    .a({\t/a/ID_rs2$0$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_2 }),
    .b({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$16$ [14],\t/a/regfile/regfile$16$ [25]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [14],\t/a/regfile/regfile$17$ [25]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1608_o,_al_u1356_o}),
    .q({\t/a/regfile/regfile$17$ [14],\t/a/regfile/regfile$17$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000000011011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b560|t/a/regfile/reg0_b568  (
    .a({\t/a/ID_rs2$0$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_2 }),
    .b({\t/a/regfile/regfile$16$ [16],\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$17$ [16],\t/a/regfile/regfile$16$ [24]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/regfile/regfile$17$ [24]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1566_o,_al_u1377_o}),
    .q({\t/a/regfile/regfile$17$ [16],\t/a/regfile/regfile$17$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b562|t/a/regfile/reg0_b566  (
    .a({\t/a/regfile/regfile$16$ [18],\t/a/ID_rs2$0$_placeOpt_7 }),
    .b({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({\t/a/ID_rs2$0$_placeOpt_7 ,\t/a/regfile/regfile$16$ [22]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [18],\t/a/regfile/regfile$17$ [22]}),
    .mi({\t/a/reg_writedat [18],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1524_o,_al_u1419_o}),
    .q({\t/a/regfile/regfile$17$ [18],\t/a/regfile/regfile$17$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b563|t/a/regfile/reg0_b564  (
    .a({\t/a/ID_rs2$0$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_1 }),
    .b({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({\t/a/regfile/regfile$16$ [19],\t/a/regfile/regfile$16$ [20]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [19],\t/a/regfile/regfile$17$ [20]}),
    .mi({\t/a/reg_writedat [19],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1503_o,_al_u1461_o}),
    .q({\t/a/regfile/regfile$17$ [19],\t/a/regfile/regfile$17$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~0*~D*C*~B*A)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~1*~D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000000100000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b576|t/a/regfile/reg0_b607  (
    .a({_al_u256_o,\t/a/ID_rs1$0$_placeOpt_10 }),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$18$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$19$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b576_sel_is_3_o ,_al_u488_o}),
    .q({\t/a/regfile/regfile$18$ [0],\t/a/regfile/regfile$18$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~B*A*~C*~D+B*A*~C*~D+~B*A*~C*D+B*A*~C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~B*A*~C*~D+B*A*~C*~D+~B*A*C*~D+B*A*C*~D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000101000001010),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b577|t/a/regfile/reg0_b592  (
    .a({\t/a/ID_rs1$1$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_2 }),
    .b({open_n38454,\t/a/ID_rs1$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$18$ [1],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [1],\t/a/regfile/regfile$18$ [16]}),
    .e({\t/a/ID_rs1$0$_placeOpt_2 ,\t/a/regfile/regfile$19$ [16]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u767_o,_al_u845_o}),
    .q({\t/a/regfile/regfile$18$ [1],\t/a/regfile/regfile$18$ [16]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b578|t/a/regfile/reg0_b606  (
    .a({\t/a/ID_rs1$0$_placeOpt_19 ,\t/a/ID_rs1$0$_placeOpt_19 }),
    .b({\t/a/ID_rs1$1$_placeOpt_19 ,\t/a/ID_rs1$1$_placeOpt_19 }),
    .c({\t/a/regfile/regfile$18$ [2],\t/a/regfile/regfile$18$ [30]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [2],\t/a/regfile/regfile$19$ [30]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u536_o,_al_u515_o}),
    .q({\t/a/regfile/regfile$18$ [2],\t/a/regfile/regfile$18$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b579|t/a/regfile/reg0_b604  (
    .a({\t/a/regfile/regfile$19$ [3],\t/a/ID_rs1$0$_placeOpt_7 }),
    .b({\t/a/regfile/regfile$18$ [3],\t/a/ID_rs1$1$_placeOpt_7 }),
    .c({\t/a/ID_rs1$0$_placeOpt_7 ,\t/a/regfile/regfile$18$ [28]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_7 ,\t/a/regfile/regfile$19$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u473_o,_al_u578_o}),
    .q({\t/a/regfile/regfile$18$ [3],\t/a/regfile/regfile$18$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1101111110001111),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b580|t/a/regfile/reg0_b605  (
    .a({\t/a/ID_rs1$0$_placeOpt_5 ,\t/a/ID_rs1$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$19$ [4],\t/a/ID_rs1$1$_placeOpt_5 }),
    .c({\t/a/ID_rs1$1$_placeOpt_5 ,\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [4],\t/a/regfile/regfile$18$ [29]}),
    .e({\t/a/ID_rs1 [2],\t/a/regfile/regfile$19$ [29]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u446_o,_al_u551_o}),
    .q({\t/a/regfile/regfile$18$ [4],\t/a/regfile/regfile$18$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b581|t/a/regfile/reg0_b602  (
    .a({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$18$ [5],\t/a/regfile/regfile$18$ [26]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [5],\t/a/regfile/regfile$19$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u431_o,_al_u620_o}),
    .q({\t/a/regfile/regfile$18$ [5],\t/a/regfile/regfile$18$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b582|t/a/regfile/reg0_b601  (
    .a({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$18$ [6],\t/a/regfile/regfile$18$ [25]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [6],\t/a/regfile/regfile$19$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u410_o,_al_u641_o}),
    .q({\t/a/regfile/regfile$18$ [6],\t/a/regfile/regfile$18$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~C*~B*~A*~D+C*~B*~A*~D+~C*B*~A*~D+C*B*~A*~D+C*B*A*~D+~C*~B*~A*D+C*~B*~A*D+~C*B*~A*D+C*B*~A*D+~C*~B*A*D+~C*B*A*D+C*B*A*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1101111111010101),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b583|t/a/regfile/reg0_b603  (
    .a({\t/a/ID_rs1$1$_placeOpt_7 ,\t/a/ID_rs1$0$_placeOpt_7 }),
    .b({\t/a/regfile/regfile$19$ [7],\t/a/ID_rs1$1$_placeOpt_7 }),
    .c({\t/a/ID_rs1$0$_placeOpt_7 ,\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [7],\t/a/regfile/regfile$18$ [27]}),
    .e({\t/a/ID_rs1 [2],\t/a/regfile/regfile$19$ [27]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u383_o,_al_u593_o}),
    .q({\t/a/regfile/regfile$18$ [7],\t/a/regfile/regfile$18$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b584|t/a/regfile/reg0_b600  (
    .a({\t/a/regfile/regfile$18$ [8],\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/regfile/regfile$19$ [8],\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/regfile/regfile$18$ [24]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/regfile/regfile$19$ [24]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u368_o,_al_u662_o}),
    .q({\t/a/regfile/regfile$18$ [8],\t/a/regfile/regfile$18$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b585|t/a/regfile/reg0_b598  (
    .a({\t/a/ID_rs1$0$_placeOpt_8 ,\t/a/ID_rs1$0$_placeOpt_8 }),
    .b({\t/a/ID_rs1$1$_placeOpt_8 ,\t/a/ID_rs1$1$_placeOpt_8 }),
    .c({\t/a/regfile/regfile$19$ [9],\t/a/ID_rs1$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [9],\t/a/regfile/regfile$18$ [22]}),
    .e({\t/a/ID_rs1$2$_placeOpt_2 ,\t/a/regfile/regfile$19$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u341_o,_al_u698_o}),
    .q({\t/a/regfile/regfile$18$ [9],\t/a/regfile/regfile$18$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b586|t/a/regfile/reg0_b599  (
    .a({\t/a/regfile/regfile$19$ [10],\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/regfile/regfile$18$ [10],\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/regfile/regfile$18$ [23]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/regfile/regfile$19$ [23]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u977_o,_al_u683_o}),
    .q({\t/a/regfile/regfile$18$ [10],\t/a/regfile/regfile$18$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b587|t/a/regfile/reg0_b596  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$19$ [11],\t/a/ID_rs1$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [11],\t/a/regfile/regfile$18$ [20]}),
    .e({\t/a/ID_rs1$2$_placeOpt_2 ,\t/a/regfile/regfile$19$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u950_o,_al_u740_o}),
    .q({\t/a/regfile/regfile$18$ [11],\t/a/regfile/regfile$18$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b588|t/a/regfile/reg0_b597  (
    .a({\t/a/regfile/regfile$19$ [12],\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/regfile/regfile$18$ [12],\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/regfile/regfile$18$ [21]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/regfile/regfile$19$ [21]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u935_o,_al_u725_o}),
    .q({\t/a/regfile/regfile$18$ [12],\t/a/regfile/regfile$18$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b589|t/a/regfile/reg0_b594  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$19$ [13],\t/a/ID_rs1$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [13],\t/a/regfile/regfile$18$ [18]}),
    .e({\t/a/ID_rs1$2$_placeOpt_2 ,\t/a/regfile/regfile$19$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u908_o,_al_u803_o}),
    .q({\t/a/regfile/regfile$18$ [13],\t/a/regfile/regfile$18$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b590|t/a/regfile/reg0_b595  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$18$ [14],\t/a/regfile/regfile$18$ [19]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [14],\t/a/regfile/regfile$19$ [19]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u893_o,_al_u788_o}),
    .q({\t/a/regfile/regfile$18$ [14],\t/a/regfile/regfile$18$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b591|t/a/regfile/reg0_b593  (
    .a({\t/a/regfile/regfile$18$ [15],\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/regfile/regfile$19$ [15],\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/regfile/regfile$18$ [17]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/regfile/regfile$19$ [17]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u872_o,_al_u830_o}),
    .q({\t/a/regfile/regfile$18$ [15],\t/a/regfile/regfile$18$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~0*~D*C*A*B)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~1*~D*C*A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b608|t/a/regfile/reg0_b638  (
    .a({\t/a/WB_rd [0],\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({_al_u256_o,\t/a/ID_rs2$1$_placeOpt_12 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2$2$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$18$ [30]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$19$ [30]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b608_sel_is_3_o ,_al_u1225_o}),
    .q({\t/a/regfile/regfile$19$ [0],\t/a/regfile/regfile$19$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b609|t/a/regfile/reg0_b639  (
    .a({\t/a/regfile/regfile$19$ [1],\t/a/ID_rs2 [0]}),
    .b({\t/a/regfile/regfile$18$ [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [1],\t/a/regfile/regfile$18$ [31]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [0],\t/a/regfile/regfile$19$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1483_o,_al_u1210_o}),
    .q({\t/a/regfile/regfile$19$ [1],\t/a/regfile/regfile$19$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b610|t/a/regfile/reg0_b637  (
    .a({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_4 }),
    .b({\t/a/ID_rs2$1$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$18$ [2],\t/a/regfile/regfile$18$ [29]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [2],\t/a/regfile/regfile$19$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1252_o,_al_u1273_o}),
    .q({\t/a/regfile/regfile$19$ [2],\t/a/regfile/regfile$19$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b611|t/a/regfile/reg0_b636  (
    .a({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/ID_rs2$1$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$19$ [3],\t/a/ID_rs2$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [3],\t/a/regfile/regfile$18$ [28]}),
    .e({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/regfile/regfile$19$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1183_o,_al_u1288_o}),
    .q({\t/a/regfile/regfile$19$ [3],\t/a/regfile/regfile$19$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000110001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b612|t/a/regfile/reg0_b635  (
    .a({\t/a/regfile/regfile$18$ [4],\t/a/ID_rs2$0$_placeOpt_4 }),
    .b({\t/a/ID_rs2$1$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$19$ [4],\t/a/regfile/regfile$18$ [27]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/regfile/regfile$19$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1168_o,_al_u1315_o}),
    .q({\t/a/regfile/regfile$19$ [4],\t/a/regfile/regfile$19$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b613|t/a/regfile/reg0_b633  (
    .a({\t/a/ID_rs2$0$_placeOpt_6 ,\t/a/ID_rs2$0$_placeOpt_6 }),
    .b({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$19$ [5],\t/a/regfile/regfile$18$ [25]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [5],\t/a/regfile/regfile$19$ [25]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1147_o,_al_u1357_o}),
    .q({\t/a/regfile/regfile$19$ [5],\t/a/regfile/regfile$19$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b614|t/a/regfile/reg0_b632  (
    .a({\t/a/ID_rs2$0$_placeOpt_6 ,\t/a/ID_rs2$0$_placeOpt_6 }),
    .b({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$18$ [6],\t/a/regfile/regfile$18$ [24]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [6],\t/a/regfile/regfile$19$ [24]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1126_o,_al_u1378_o}),
    .q({\t/a/regfile/regfile$19$ [6],\t/a/regfile/regfile$19$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0001000010110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b615|t/a/regfile/reg0_b630  (
    .a({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$18$ [7],\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/regfile/regfile$18$ [22]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [7],\t/a/regfile/regfile$19$ [22]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1105_o,_al_u1420_o}),
    .q({\t/a/regfile/regfile$19$ [7],\t/a/regfile/regfile$19$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b616|t/a/regfile/reg0_b634  (
    .a({\t/a/ID_rs2$0$_placeOpt_6 ,\t/a/ID_rs2$0$_placeOpt_6 }),
    .b({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$19$ [8],\t/a/ID_rs2$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [8],\t/a/regfile/regfile$18$ [26]}),
    .e({\t/a/ID_rs2$2$_placeOpt_9 ,\t/a/regfile/regfile$19$ [26]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1078_o,_al_u1330_o}),
    .q({\t/a/regfile/regfile$19$ [8],\t/a/regfile/regfile$19$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b617|t/a/regfile/reg0_b628  (
    .a({\t/a/regfile/regfile$18$ [9],\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$19$ [9],\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/regfile/regfile$18$ [20]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/regfile/regfile$19$ [20]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1063_o,_al_u1462_o}),
    .q({\t/a/regfile/regfile$19$ [9],\t/a/regfile/regfile$19$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b618|t/a/regfile/reg0_b631  (
    .a({\t/a/ID_rs2$0$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_2 }),
    .b({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$19$ [10],\t/a/ID_rs2$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [10],\t/a/regfile/regfile$18$ [23]}),
    .e({\t/a/ID_rs2$2$_placeOpt_9 ,\t/a/regfile/regfile$19$ [23]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1687_o,_al_u1393_o}),
    .q({\t/a/regfile/regfile$19$ [10],\t/a/regfile/regfile$19$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b619|t/a/regfile/reg0_b627  (
    .a({\t/a/regfile/regfile$18$ [11],\t/a/ID_rs2$0$_placeOpt_7 }),
    .b({\t/a/regfile/regfile$19$ [11],\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({\t/a/ID_rs2$0$_placeOpt_7 ,\t/a/regfile/regfile$18$ [19]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/regfile/regfile$19$ [19]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1672_o,_al_u1504_o}),
    .q({\t/a/regfile/regfile$19$ [11],\t/a/regfile/regfile$19$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b620|t/a/regfile/reg0_b629  (
    .a({\t/a/ID_rs2$0$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_2 }),
    .b({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$19$ [12],\t/a/ID_rs2$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [12],\t/a/regfile/regfile$18$ [21]}),
    .e({\t/a/ID_rs2$2$_placeOpt_9 ,\t/a/regfile/regfile$19$ [21]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1645_o,_al_u1435_o}),
    .q({\t/a/regfile/regfile$19$ [12],\t/a/regfile/regfile$19$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b621|t/a/regfile/reg0_b626  (
    .a({\t/a/regfile/regfile$18$ [13],\t/a/ID_rs2$0$_placeOpt_7 }),
    .b({\t/a/regfile/regfile$19$ [13],\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({\t/a/ID_rs2$0$_placeOpt_7 ,\t/a/regfile/regfile$18$ [18]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/regfile/regfile$19$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1630_o,_al_u1525_o}),
    .q({\t/a/regfile/regfile$19$ [13],\t/a/regfile/regfile$19$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b622|t/a/regfile/reg0_b624  (
    .a({\t/a/ID_rs2$0$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_1 }),
    .b({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({\t/a/regfile/regfile$19$ [14],\t/a/regfile/regfile$18$ [16]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [14],\t/a/regfile/regfile$19$ [16]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1609_o,_al_u1567_o}),
    .q({\t/a/regfile/regfile$19$ [14],\t/a/regfile/regfile$19$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b623|t/a/regfile/reg0_b625  (
    .a({\t/a/ID_rs2$0$_placeOpt_6 ,\t/a/ID_rs2$0$_placeOpt_6 }),
    .b({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$19$ [15],\t/a/ID_rs2$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [15],\t/a/regfile/regfile$18$ [17]}),
    .e({\t/a/ID_rs2$2$_placeOpt_2 ,\t/a/regfile/regfile$19$ [17]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1582_o,_al_u1540_o}),
    .q({\t/a/regfile/regfile$19$ [15],\t/a/regfile/regfile$19$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b641|t/a/regfile/reg0_b670  (
    .a({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/ID_rs1$0$_placeOpt_13 }),
    .b({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/ID_rs1$1$_placeOpt_13 }),
    .c({\t/a/regfile/regfile$20$ [1],\t/a/regfile/regfile$20$ [30]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [1],\t/a/regfile/regfile$21$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u764_o,_al_u512_o}),
    .q({\t/a/regfile/regfile$20$ [1],\t/a/regfile/regfile$20$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b642|t/a/regfile/reg0_b668  (
    .a({\t/a/ID_rs1$0$_placeOpt_5 ,\t/a/ID_rs1$0$_placeOpt_5 }),
    .b({\t/a/ID_rs1$1$_placeOpt_5 ,\t/a/ID_rs1$1$_placeOpt_5 }),
    .c({\t/a/regfile/regfile$21$ [2],\t/a/regfile/regfile$20$ [28]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$20$ [2],\t/a/regfile/regfile$21$ [28]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u533_o,_al_u575_o}),
    .q({\t/a/regfile/regfile$20$ [2],\t/a/regfile/regfile$20$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b643|t/a/regfile/reg0_b666  (
    .a({\t/a/regfile/regfile$21$ [3],\t/a/ID_rs1 [0]}),
    .b({\t/a/regfile/regfile$20$ [3],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [1],\t/a/regfile/regfile$20$ [26]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [0],\t/a/regfile/regfile$21$ [26]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u470_o,_al_u617_o}),
    .q({\t/a/regfile/regfile$20$ [3],\t/a/regfile/regfile$20$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b645|t/a/regfile/reg0_b665  (
    .a({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$20$ [5],\t/a/regfile/regfile$20$ [25]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [5],\t/a/regfile/regfile$21$ [25]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u428_o,_al_u638_o}),
    .q({\t/a/regfile/regfile$20$ [5],\t/a/regfile/regfile$20$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b646|t/a/regfile/reg0_b664  (
    .a({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$21$ [6],\t/a/regfile/regfile$20$ [24]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$20$ [6],\t/a/regfile/regfile$21$ [24]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u407_o,_al_u659_o}),
    .q({\t/a/regfile/regfile$20$ [6],\t/a/regfile/regfile$20$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b648|t/a/regfile/reg0_b663  (
    .a({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/regfile/regfile$20$ [8],\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/regfile/regfile$20$ [23]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [8],\t/a/regfile/regfile$21$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u365_o,_al_u680_o}),
    .q({\t/a/regfile/regfile$20$ [8],\t/a/regfile/regfile$20$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b650|t/a/regfile/reg0_b661  (
    .a({\t/a/regfile/regfile$21$ [10],\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/regfile/regfile$20$ [10],\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/regfile/regfile$20$ [21]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/regfile/regfile$21$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u974_o,_al_u722_o}),
    .q({\t/a/regfile/regfile$20$ [10],\t/a/regfile/regfile$20$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b652|t/a/regfile/reg0_b659  (
    .a({\t/a/regfile/regfile$20$ [12],\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/regfile/regfile$20$ [19]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [12],\t/a/regfile/regfile$21$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u932_o,_al_u785_o}),
    .q({\t/a/regfile/regfile$20$ [12],\t/a/regfile/regfile$20$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b654|t/a/regfile/reg0_b657  (
    .a({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/regfile/regfile$20$ [14],\t/a/regfile/regfile$20$ [17]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [14],\t/a/regfile/regfile$21$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u890_o,_al_u827_o}),
    .q({\t/a/regfile/regfile$20$ [14],\t/a/regfile/regfile$20$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b65|t/a/regfile/reg0_b68  (
    .a({\t/a/ID_rs1$0$_placeOpt_16 ,\t/a/ID_rs1$0$_placeOpt_16 }),
    .b({\t/a/ID_rs1$1$_placeOpt_10 ,\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/regfile/regfile$3$ [1],\t/a/regfile/regfile$3$ [4]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [1],\t/a/regfile/regfile$2$ [4]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u757_o,_al_u452_o}),
    .q({\t/a/regfile/regfile$2$ [1],\t/a/regfile/regfile$2$ [4]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b66|t/a/regfile/reg0_b67  (
    .a({\t/a/ID_rs1$0$_placeOpt_10 ,\t/a/ID_rs1$0$_placeOpt_10 }),
    .b({\t/a/ID_rs1$1$_placeOpt_10 ,\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/regfile/regfile$2$ [2],\t/a/regfile/regfile$2$ [3]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$3$ [2],\t/a/regfile/regfile$3$ [3]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u526_o,_al_u463_o}),
    .q({\t/a/regfile/regfile$2$ [2],\t/a/regfile/regfile$2$ [3]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b673|t/a/regfile/reg0_b703  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$20$ [1],\t/a/regfile/regfile$20$ [31]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [1],\t/a/regfile/regfile$21$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1480_o,_al_u1207_o}),
    .q({\t/a/regfile/regfile$21$ [1],\t/a/regfile/regfile$21$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b674|t/a/regfile/reg0_b701  (
    .a({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_4 }),
    .b({\t/a/ID_rs2$1$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$20$ [2],\t/a/regfile/regfile$20$ [29]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [2],\t/a/regfile/regfile$21$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1249_o,_al_u1270_o}),
    .q({\t/a/regfile/regfile$21$ [2],\t/a/regfile/regfile$21$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b676|t/a/regfile/reg0_b699  (
    .a({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_4 }),
    .b({\t/a/regfile/regfile$20$ [4],\t/a/ID_rs2$1$_placeOpt_1 }),
    .c({\t/a/ID_rs2$1$_placeOpt_1 ,\t/a/regfile/regfile$20$ [27]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [4],\t/a/regfile/regfile$21$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1165_o,_al_u1312_o}),
    .q({\t/a/regfile/regfile$21$ [4],\t/a/regfile/regfile$21$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b677|t/a/regfile/reg0_b697  (
    .a({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs2$0$_placeOpt_12 }),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_5 }),
    .c({\t/a/regfile/regfile$21$ [5],\t/a/regfile/regfile$20$ [25]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$20$ [5],\t/a/regfile/regfile$21$ [25]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1144_o,_al_u1354_o}),
    .q({\t/a/regfile/regfile$21$ [5],\t/a/regfile/regfile$21$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b678|t/a/regfile/reg0_b696  (
    .a({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs2$0$_placeOpt_12 }),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_5 }),
    .c({\t/a/regfile/regfile$20$ [6],\t/a/regfile/regfile$20$ [24]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [6],\t/a/regfile/regfile$21$ [24]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1123_o,_al_u1375_o}),
    .q({\t/a/regfile/regfile$21$ [6],\t/a/regfile/regfile$21$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b679|t/a/regfile/reg0_b694  (
    .a({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$20$ [7],\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/regfile/regfile$20$ [22]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [7],\t/a/regfile/regfile$21$ [22]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1102_o,_al_u1417_o}),
    .q({\t/a/regfile/regfile$21$ [7],\t/a/regfile/regfile$21$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b681|t/a/regfile/reg0_b692  (
    .a({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$20$ [9],\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/regfile/regfile$20$ [20]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [9],\t/a/regfile/regfile$21$ [20]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1060_o,_al_u1459_o}),
    .q({\t/a/regfile/regfile$21$ [9],\t/a/regfile/regfile$21$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b683|t/a/regfile/reg0_b691  (
    .a({\t/a/regfile/regfile$21$ [11],\t/a/ID_rs2$0$_placeOpt_8 }),
    .b({\t/a/regfile/regfile$20$ [11],\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/regfile/regfile$20$ [19]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_8 ,\t/a/regfile/regfile$21$ [19]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1669_o,_al_u1501_o}),
    .q({\t/a/regfile/regfile$21$ [11],\t/a/regfile/regfile$21$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b685|t/a/regfile/reg0_b690  (
    .a({\t/a/regfile/regfile$21$ [13],\t/a/ID_rs2$0$_placeOpt_7 }),
    .b({\t/a/regfile/regfile$20$ [13],\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/regfile/regfile$20$ [18]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_7 ,\t/a/regfile/regfile$21$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1627_o,_al_u1522_o}),
    .q({\t/a/regfile/regfile$21$ [13],\t/a/regfile/regfile$21$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b686|t/a/regfile/reg0_b688  (
    .a({\t/a/ID_rs2$0$_placeOpt_8 ,\t/a/ID_rs2$0$_placeOpt_8 }),
    .b({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$20$ [14],\t/a/regfile/regfile$20$ [16]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [14],\t/a/regfile/regfile$21$ [16]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1606_o,_al_u1564_o}),
    .q({\t/a/regfile/regfile$21$ [14],\t/a/regfile/regfile$21$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~0*D*C*~B*A)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~1*D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b704|t/a/regfile/reg0_b735  (
    .a({_al_u256_o,\t/a/ID_rs1$0$_placeOpt_10 }),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1$2$_placeOpt_4 }),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$22$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$23$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b704_sel_is_3_o ,_al_u486_o}),
    .q({\t/a/regfile/regfile$22$ [0],\t/a/regfile/regfile$22$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*D*~C*~B+A*D*~C*~B+A*D*C*~B+~A*D*~C*B+A*D*~C*B+A*D*C*B"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*D*~C*~B+~A*D*~C*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b1010111100000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0000010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b705|t/a/regfile/reg0_b720  (
    .a({\t/a/ID_rs1$0$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_2 }),
    .b({open_n39170,\t/a/ID_rs1$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$22$ [1],\t/a/ID_rs1$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_2 ,\t/a/regfile/regfile$22$ [16]}),
    .e({\t/a/regfile/regfile$23$ [1],\t/a/regfile/regfile$23$ [16]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u765_o,_al_u843_o}),
    .q({\t/a/regfile/regfile$22$ [1],\t/a/regfile/regfile$22$ [16]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b706|t/a/regfile/reg0_b734  (
    .a({\t/a/ID_rs1$0$_placeOpt_19 ,\t/a/ID_rs1$0$_placeOpt_19 }),
    .b({\t/a/ID_rs1$1$_placeOpt_19 ,\t/a/ID_rs1$1$_placeOpt_19 }),
    .c({\t/a/regfile/regfile$23$ [2],\t/a/regfile/regfile$22$ [30]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [2],\t/a/regfile/regfile$23$ [30]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u534_o,_al_u513_o}),
    .q({\t/a/regfile/regfile$22$ [2],\t/a/regfile/regfile$22$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b707|t/a/regfile/reg0_b732  (
    .a({\t/a/regfile/regfile$23$ [3],\t/a/ID_rs1$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$22$ [3],\t/a/ID_rs1$1$_placeOpt_5 }),
    .c({\t/a/ID_rs1$1$_placeOpt_5 ,\t/a/regfile/regfile$22$ [28]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_5 ,\t/a/regfile/regfile$23$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u471_o,_al_u576_o}),
    .q({\t/a/regfile/regfile$22$ [3],\t/a/regfile/regfile$22$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1101111110001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b708|t/a/regfile/reg0_b733  (
    .a({\t/a/ID_rs1$0$_placeOpt_5 ,\t/a/ID_rs1$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$23$ [4],\t/a/ID_rs1$1$_placeOpt_5 }),
    .c({\t/a/ID_rs1$1$_placeOpt_5 ,\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [4],\t/a/regfile/regfile$22$ [29]}),
    .e({\t/a/ID_rs1 [2],\t/a/regfile/regfile$23$ [29]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u444_o,_al_u549_o}),
    .q({\t/a/regfile/regfile$22$ [4],\t/a/regfile/regfile$22$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b709|t/a/regfile/reg0_b730  (
    .a({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$22$ [5],\t/a/regfile/regfile$22$ [26]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [5],\t/a/regfile/regfile$23$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u429_o,_al_u618_o}),
    .q({\t/a/regfile/regfile$22$ [5],\t/a/regfile/regfile$22$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b710|t/a/regfile/reg0_b729  (
    .a({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$22$ [6],\t/a/regfile/regfile$22$ [25]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [6],\t/a/regfile/regfile$23$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u408_o,_al_u639_o}),
    .q({\t/a/regfile/regfile$22$ [6],\t/a/regfile/regfile$22$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1011111110110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b711|t/a/regfile/reg0_b731  (
    .a({\t/a/regfile/regfile$23$ [7],\t/a/ID_rs1$0$_placeOpt_5 }),
    .b({\t/a/ID_rs1$1$_placeOpt_5 ,\t/a/ID_rs1$1$_placeOpt_5 }),
    .c({\t/a/ID_rs1$0$_placeOpt_5 ,\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [7],\t/a/regfile/regfile$22$ [27]}),
    .e({\t/a/ID_rs1 [2],\t/a/regfile/regfile$23$ [27]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u381_o,_al_u591_o}),
    .q({\t/a/regfile/regfile$22$ [7],\t/a/regfile/regfile$22$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b712|t/a/regfile/reg0_b728  (
    .a({\t/a/regfile/regfile$23$ [8],\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/regfile/regfile$22$ [8],\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/regfile/regfile$22$ [24]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/regfile/regfile$23$ [24]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u366_o,_al_u660_o}),
    .q({\t/a/regfile/regfile$22$ [8],\t/a/regfile/regfile$22$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111011110110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b713|t/a/regfile/reg0_b726  (
    .a({\t/a/ID_rs1$0$_placeOpt_7 ,\t/a/ID_rs1$0$_placeOpt_7 }),
    .b({\t/a/ID_rs1$1$_placeOpt_7 ,\t/a/ID_rs1$1$_placeOpt_7 }),
    .c({\t/a/regfile/regfile$23$ [9],\t/a/ID_rs1$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [9],\t/a/regfile/regfile$22$ [22]}),
    .e({\t/a/ID_rs1$2$_placeOpt_2 ,\t/a/regfile/regfile$23$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u339_o,_al_u696_o}),
    .q({\t/a/regfile/regfile$22$ [9],\t/a/regfile/regfile$22$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b714|t/a/regfile/reg0_b727  (
    .a({\t/a/regfile/regfile$23$ [10],\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/regfile/regfile$22$ [10],\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/regfile/regfile$22$ [23]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/regfile/regfile$23$ [23]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u975_o,_al_u681_o}),
    .q({\t/a/regfile/regfile$22$ [10],\t/a/regfile/regfile$22$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111001110111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b715|t/a/regfile/reg0_b724  (
    .a({\t/a/regfile/regfile$22$ [11],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$23$ [11],\t/a/ID_rs1$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [0],\t/a/regfile/regfile$22$ [20]}),
    .e({\t/a/ID_rs1$2$_placeOpt_2 ,\t/a/regfile/regfile$23$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u948_o,_al_u738_o}),
    .q({\t/a/regfile/regfile$22$ [11],\t/a/regfile/regfile$22$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b716|t/a/regfile/reg0_b725  (
    .a({\t/a/regfile/regfile$22$ [12],\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/regfile/regfile$23$ [12],\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/regfile/regfile$22$ [21]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/regfile/regfile$23$ [21]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u933_o,_al_u723_o}),
    .q({\t/a/regfile/regfile$22$ [12],\t/a/regfile/regfile$22$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111011110110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b717|t/a/regfile/reg0_b722  (
    .a({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/regfile/regfile$23$ [13],\t/a/ID_rs1$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [13],\t/a/regfile/regfile$22$ [18]}),
    .e({\t/a/ID_rs1$2$_placeOpt_7 ,\t/a/regfile/regfile$23$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u906_o,_al_u801_o}),
    .q({\t/a/regfile/regfile$22$ [13],\t/a/regfile/regfile$22$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b718|t/a/regfile/reg0_b723  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$22$ [14],\t/a/regfile/regfile$22$ [19]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [14],\t/a/regfile/regfile$23$ [19]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u891_o,_al_u786_o}),
    .q({\t/a/regfile/regfile$22$ [14],\t/a/regfile/regfile$22$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b719|t/a/regfile/reg0_b721  (
    .a({\t/a/regfile/regfile$22$ [15],\t/a/ID_rs1$0$_placeOpt_4 }),
    .b({\t/a/regfile/regfile$23$ [15],\t/a/ID_rs1$1$_placeOpt_4 }),
    .c({\t/a/ID_rs1$0$_placeOpt_4 ,\t/a/regfile/regfile$22$ [17]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_4 ,\t/a/regfile/regfile$23$ [17]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u870_o,_al_u828_o}),
    .q({\t/a/regfile/regfile$22$ [15],\t/a/regfile/regfile$22$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~0*D*C*B*A)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~1*D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b736|t/a/regfile/reg0_b766  (
    .a({_al_u256_o,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2$1$_placeOpt_11 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2$2$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$22$ [30]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$23$ [30]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b736_sel_is_3_o ,_al_u1223_o}),
    .q({\t/a/regfile/regfile$23$ [0],\t/a/regfile/regfile$23$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b737|t/a/regfile/reg0_b767  (
    .a({\t/a/regfile/regfile$23$ [1],\t/a/ID_rs2 [0]}),
    .b({\t/a/regfile/regfile$22$ [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [1],\t/a/regfile/regfile$22$ [31]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [0],\t/a/regfile/regfile$23$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1481_o,_al_u1208_o}),
    .q({\t/a/regfile/regfile$23$ [1],\t/a/regfile/regfile$23$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b738|t/a/regfile/reg0_b765  (
    .a({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_4 }),
    .b({\t/a/ID_rs2$1$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$22$ [2],\t/a/regfile/regfile$22$ [29]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [2],\t/a/regfile/regfile$23$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1250_o,_al_u1271_o}),
    .q({\t/a/regfile/regfile$23$ [2],\t/a/regfile/regfile$23$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111011110110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b739|t/a/regfile/reg0_b764  (
    .a({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_4 }),
    .b({\t/a/ID_rs2$1$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$23$ [3],\t/a/ID_rs2$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [3],\t/a/regfile/regfile$22$ [28]}),
    .e({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/regfile/regfile$23$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1181_o,_al_u1286_o}),
    .q({\t/a/regfile/regfile$23$ [3],\t/a/regfile/regfile$23$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(A*~(C)*~(D)+A*C*~(D)+~(A)*C*D+A*C*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000110001000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b740|t/a/regfile/reg0_b763  (
    .a({\t/a/regfile/regfile$22$ [4],\t/a/ID_rs2$0$_placeOpt_4 }),
    .b({\t/a/ID_rs2$1$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$23$ [4],\t/a/regfile/regfile$22$ [27]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/regfile/regfile$23$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1166_o,_al_u1313_o}),
    .q({\t/a/regfile/regfile$23$ [4],\t/a/regfile/regfile$23$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b741|t/a/regfile/reg0_b761  (
    .a({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs2$0$_placeOpt_12 }),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_5 }),
    .c({\t/a/regfile/regfile$22$ [5],\t/a/regfile/regfile$22$ [25]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [5],\t/a/regfile/regfile$23$ [25]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1145_o,_al_u1355_o}),
    .q({\t/a/regfile/regfile$23$ [5],\t/a/regfile/regfile$23$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b742|t/a/regfile/reg0_b760  (
    .a({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs2$0$_placeOpt_12 }),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_5 }),
    .c({\t/a/regfile/regfile$22$ [6],\t/a/regfile/regfile$22$ [24]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [6],\t/a/regfile/regfile$23$ [24]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1124_o,_al_u1376_o}),
    .q({\t/a/regfile/regfile$23$ [6],\t/a/regfile/regfile$23$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0001101100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b743|t/a/regfile/reg0_b758  (
    .a({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$22$ [7],\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/regfile/regfile$23$ [7],\t/a/regfile/regfile$22$ [22]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/regfile/regfile$23$ [22]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1103_o,_al_u1418_o}),
    .q({\t/a/regfile/regfile$23$ [7],\t/a/regfile/regfile$23$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111011110110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b744|t/a/regfile/reg0_b762  (
    .a({\t/a/ID_rs2$0$_placeOpt_6 ,\t/a/ID_rs2$0$_placeOpt_6 }),
    .b({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$23$ [8],\t/a/ID_rs2$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [8],\t/a/regfile/regfile$22$ [26]}),
    .e({\t/a/ID_rs2$2$_placeOpt_9 ,\t/a/regfile/regfile$23$ [26]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1076_o,_al_u1328_o}),
    .q({\t/a/regfile/regfile$23$ [8],\t/a/regfile/regfile$23$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b745|t/a/regfile/reg0_b756  (
    .a({\t/a/regfile/regfile$22$ [9],\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$23$ [9],\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/regfile/regfile$22$ [20]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/regfile/regfile$23$ [20]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1061_o,_al_u1460_o}),
    .q({\t/a/regfile/regfile$23$ [9],\t/a/regfile/regfile$23$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111011110110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b746|t/a/regfile/reg0_b759  (
    .a({\t/a/ID_rs2$0$_placeOpt_6 ,\t/a/ID_rs2$0$_placeOpt_6 }),
    .b({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$23$ [10],\t/a/ID_rs2$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [10],\t/a/regfile/regfile$22$ [23]}),
    .e({\t/a/ID_rs2$2$_placeOpt_9 ,\t/a/regfile/regfile$23$ [23]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1685_o,_al_u1391_o}),
    .q({\t/a/regfile/regfile$23$ [10],\t/a/regfile/regfile$23$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0100010000001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b747|t/a/regfile/reg0_b755  (
    .a({\t/a/regfile/regfile$23$ [11],\t/a/ID_rs2$0$_placeOpt_1 }),
    .b({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({\t/a/regfile/regfile$22$ [11],\t/a/regfile/regfile$22$ [19]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_1 ,\t/a/regfile/regfile$23$ [19]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1670_o,_al_u1502_o}),
    .q({\t/a/regfile/regfile$23$ [11],\t/a/regfile/regfile$23$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111011110110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b748|t/a/regfile/reg0_b757  (
    .a({\t/a/ID_rs2$0$_placeOpt_6 ,\t/a/ID_rs2$0$_placeOpt_6 }),
    .b({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/ID_rs2$1$_placeOpt_4 }),
    .c({\t/a/regfile/regfile$23$ [12],\t/a/ID_rs2$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [12],\t/a/regfile/regfile$22$ [21]}),
    .e({\t/a/ID_rs2$2$_placeOpt_9 ,\t/a/regfile/regfile$23$ [21]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1643_o,_al_u1433_o}),
    .q({\t/a/regfile/regfile$23$ [12],\t/a/regfile/regfile$23$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b749|t/a/regfile/reg0_b754  (
    .a({\t/a/regfile/regfile$22$ [13],\t/a/ID_rs2$0$_placeOpt_7 }),
    .b({\t/a/regfile/regfile$23$ [13],\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({\t/a/ID_rs2$0$_placeOpt_7 ,\t/a/regfile/regfile$22$ [18]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/regfile/regfile$23$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1628_o,_al_u1523_o}),
    .q({\t/a/regfile/regfile$23$ [13],\t/a/regfile/regfile$23$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b750|t/a/regfile/reg0_b752  (
    .a({\t/a/ID_rs2$0$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_1 }),
    .b({\t/a/ID_rs2$1$_placeOpt_16 ,\t/a/ID_rs2$1$_placeOpt_16 }),
    .c({\t/a/regfile/regfile$22$ [14],\t/a/regfile/regfile$22$ [16]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [14],\t/a/regfile/regfile$23$ [16]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1607_o,_al_u1565_o}),
    .q({\t/a/regfile/regfile$23$ [14],\t/a/regfile/regfile$23$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("0"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111011110110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b751|t/a/regfile/reg0_b753  (
    .a({\t/a/ID_rs2$0$_placeOpt_12 ,\t/a/ID_rs2$0$_placeOpt_12 }),
    .b({\t/a/ID_rs2$1$_placeOpt_5 ,\t/a/ID_rs2$1$_placeOpt_5 }),
    .c({\t/a/regfile/regfile$23$ [15],\t/a/ID_rs2$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [15],\t/a/regfile/regfile$22$ [17]}),
    .e({\t/a/ID_rs2$2$_placeOpt_2 ,\t/a/regfile/regfile$23$ [17]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1580_o,_al_u1538_o}),
    .q({\t/a/regfile/regfile$23$ [15],\t/a/regfile/regfile$23$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b768|t/a/regfile/reg0_b798  (
    .a({_al_u256_o,_al_u519_o}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1$0$_placeOpt_10 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1$1$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$24$ [30]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$25$ [30]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b768_sel_is_3_o ,_al_u520_o}),
    .q({\t/a/regfile/regfile$24$ [0],\t/a/regfile/regfile$24$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b769|t/a/regfile/reg0_b796  (
    .a({_al_u771_o,_al_u582_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_5 ,\t/a/ID_rs1$0$_placeOpt_5 }),
    .c({\t/a/ID_rs1$1$_placeOpt_5 ,\t/a/ID_rs1$1$_placeOpt_5 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [1],\t/a/regfile/regfile$24$ [28]}),
    .e({\t/a/regfile/regfile$25$ [1],\t/a/regfile/regfile$25$ [28]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u772_o,_al_u583_o}),
    .q({\t/a/regfile/regfile$24$ [1],\t/a/regfile/regfile$24$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b770|t/a/regfile/reg0_b794  (
    .a({_al_u540_o,_al_u624_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_3 ,\t/a/ID_rs1$0$_placeOpt_3 }),
    .c({\t/a/ID_rs1$1$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [2],\t/a/regfile/regfile$24$ [26]}),
    .e({\t/a/regfile/regfile$25$ [2],\t/a/regfile/regfile$25$ [26]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u541_o,_al_u625_o}),
    .q({\t/a/regfile/regfile$24$ [2],\t/a/regfile/regfile$24$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b771|t/a/regfile/reg0_b793  (
    .a({_al_u477_o,_al_u645_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_3 ,\t/a/ID_rs1$0$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$24$ [3],\t/a/ID_rs1$1$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_3 ,\t/a/regfile/regfile$24$ [25]}),
    .e({\t/a/regfile/regfile$25$ [3],\t/a/regfile/regfile$25$ [25]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u478_o,_al_u646_o}),
    .q({\t/a/regfile/regfile$24$ [3],\t/a/regfile/regfile$24$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~B*~D*~C*~A+B*~D*~C*~A+B*~D*C*~A+~B*~D*~C*A+B*~D*~C*A+B*~D*C*A"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~B*~D*~C*~A+~B*~D*~C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000011001111),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b772|t/a/regfile/reg0_b792  (
    .a({open_n39658,_al_u666_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_15 ,\t/a/ID_rs1$0$_placeOpt_15 }),
    .c({\t/a/regfile/regfile$24$ [4],\t/a/ID_rs1$1$_placeOpt_15 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_15 ,\t/a/regfile/regfile$24$ [24]}),
    .e({\t/a/regfile/regfile$25$ [4],\t/a/regfile/regfile$25$ [24]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u441_o,_al_u667_o}),
    .q({\t/a/regfile/regfile$24$ [4],\t/a/regfile/regfile$24$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b773|t/a/regfile/reg0_b791  (
    .a({_al_u435_o,_al_u687_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .c({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/ID_rs1$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [5],\t/a/regfile/regfile$24$ [23]}),
    .e({\t/a/regfile/regfile$25$ [5],\t/a/regfile/regfile$25$ [23]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u436_o,_al_u688_o}),
    .q({\t/a/regfile/regfile$24$ [5],\t/a/regfile/regfile$24$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b774|t/a/regfile/reg0_b789  (
    .a({_al_u414_o,_al_u729_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .c({\t/a/regfile/regfile$24$ [6],\t/a/ID_rs1$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/regfile/regfile$24$ [21]}),
    .e({\t/a/regfile/regfile$25$ [6],\t/a/regfile/regfile$25$ [21]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u415_o,_al_u730_o}),
    .q({\t/a/regfile/regfile$24$ [6],\t/a/regfile/regfile$24$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+A*~B*C*~D+~A*~B*~C*D+A*~B*~C*D+A*~B*C*D"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0010001100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b775|t/a/regfile/reg0_b787  (
    .a({\t/a/ID_rs1$0$_placeOpt_8 ,_al_u792_o}),
    .b({\t/a/ID_rs1$1$_placeOpt_8 ,\t/a/ID_rs1$0$_placeOpt_8 }),
    .c({\t/a/regfile/regfile$24$ [7],\t/a/ID_rs1$1$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({open_n39704,\t/a/regfile/regfile$24$ [19]}),
    .e({\t/a/regfile/regfile$25$ [7],\t/a/regfile/regfile$25$ [19]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u378_o,_al_u793_o}),
    .q({\t/a/regfile/regfile$24$ [7],\t/a/regfile/regfile$24$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b776|t/a/regfile/reg0_b785  (
    .a({_al_u372_o,_al_u834_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_3 ,\t/a/ID_rs1$0$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$24$ [8],\t/a/ID_rs1$1$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_3 ,\t/a/regfile/regfile$24$ [17]}),
    .e({\t/a/regfile/regfile$25$ [8],\t/a/regfile/regfile$25$ [17]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u373_o,_al_u835_o}),
    .q({\t/a/regfile/regfile$24$ [8],\t/a/regfile/regfile$24$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~C*~A*~D*~B+C*~A*~D*~B+C*~A*D*~B+~C*~A*~D*B+C*~A*~D*B+C*~A*D*B"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~C*~A*~D*~B+~C*~A*~D*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0101000001010101),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b777|t/a/regfile/reg0_b783  (
    .a({\t/a/ID_rs1$1$_placeOpt_8 ,_al_u876_o}),
    .b({open_n39735,\t/a/ID_rs1$0$_placeOpt_8 }),
    .c({\t/a/ID_rs1$0$_placeOpt_8 ,\t/a/ID_rs1$1$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [9],\t/a/regfile/regfile$24$ [15]}),
    .e({\t/a/regfile/regfile$25$ [9],\t/a/regfile/regfile$25$ [15]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u336_o,_al_u877_o}),
    .q({\t/a/regfile/regfile$24$ [9],\t/a/regfile/regfile$24$ [15]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b778|t/a/regfile/reg0_b782  (
    .a({_al_u981_o,_al_u897_o}),
    .b({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .c({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/ID_rs1$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [10],\t/a/regfile/regfile$24$ [14]}),
    .e({\t/a/regfile/regfile$25$ [10],\t/a/regfile/regfile$25$ [14]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u982_o,_al_u898_o}),
    .q({\t/a/regfile/regfile$24$ [10],\t/a/regfile/regfile$24$ [14]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~A*~C*~D*~B+A*~C*~D*~B+A*~C*D*~B+~A*~C*~D*B+A*~C*~D*B+A*~C*D*B"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~A*~C*~D*~B+~A*~C*~D*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000101000001111),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b779|t/a/regfile/reg0_b780  (
    .a({\t/a/ID_rs1$0$_placeOpt_3 ,_al_u939_o}),
    .b({open_n39766,\t/a/ID_rs1$0$_placeOpt_3 }),
    .c({\t/a/ID_rs1$1$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [11],\t/a/regfile/regfile$24$ [12]}),
    .e({\t/a/regfile/regfile$25$ [11],\t/a/regfile/regfile$25$ [12]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u945_o,_al_u940_o}),
    .q({\t/a/regfile/regfile$24$ [11],\t/a/regfile/regfile$24$ [12]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b781|t/a/regfile/reg0_b799  (
    .a({\t/a/ID_rs1$0$_placeOpt_19 ,\t/a/ID_rs1$0$_placeOpt_19 }),
    .b({\t/a/ID_rs1$1$_placeOpt_19 ,\t/a/ID_rs1$1$_placeOpt_19 }),
    .c({\t/a/regfile/regfile$24$ [13],\t/a/regfile/regfile$24$ [31]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [13],\t/a/regfile/regfile$25$ [31]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u903_o,_al_u483_o}),
    .q({\t/a/regfile/regfile$24$ [13],\t/a/regfile/regfile$24$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b784|t/a/regfile/reg0_b797  (
    .a({\t/a/regfile/regfile$24$ [16],\t/a/ID_rs1$0$_placeOpt_5 }),
    .b({\t/a/ID_rs1$1$_placeOpt_5 ,\t/a/ID_rs1$1$_placeOpt_5 }),
    .c({\t/a/ID_rs1$0$_placeOpt_5 ,\t/a/regfile/regfile$24$ [29]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [16],\t/a/regfile/regfile$25$ [29]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u840_o,_al_u546_o}),
    .q({\t/a/regfile/regfile$24$ [16],\t/a/regfile/regfile$24$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b786|t/a/regfile/reg0_b795  (
    .a({\t/a/ID_rs1$0$_placeOpt_8 ,\t/a/ID_rs1$0$_placeOpt_8 }),
    .b({\t/a/regfile/regfile$24$ [18],\t/a/ID_rs1$1$_placeOpt_8 }),
    .c({\t/a/ID_rs1$1$_placeOpt_8 ,\t/a/regfile/regfile$24$ [27]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [18],\t/a/regfile/regfile$25$ [27]}),
    .mi({\t/a/reg_writedat [18],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u798_o,_al_u588_o}),
    .q({\t/a/regfile/regfile$24$ [18],\t/a/regfile/regfile$24$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000000011011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b788|t/a/regfile/reg0_b790  (
    .a({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/regfile/regfile$24$ [20],\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/regfile/regfile$25$ [20],\t/a/regfile/regfile$24$ [22]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/regfile/regfile$25$ [22]}),
    .mi({\t/a/reg_writedat [20],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u735_o,_al_u693_o}),
    .q({\t/a/regfile/regfile$24$ [20],\t/a/regfile/regfile$24$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*~D*~C*A*B)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*~D*~C*A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b800|t/a/regfile/reg0_b831  (
    .a({\t/a/WB_rd [0],_al_u1214_o}),
    .b({_al_u256_o,\t/a/ID_rs2$0$_placeOpt_22 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2$1$_placeOpt_11 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$24$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$25$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b800_sel_is_3_o ,_al_u1215_o}),
    .q({\t/a/regfile/regfile$25$ [0],\t/a/regfile/regfile$25$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b801|t/a/regfile/reg0_b829  (
    .a({_al_u1487_o,_al_u1277_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_4 }),
    .c({\t/a/ID_rs2$1$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [1],\t/a/regfile/regfile$24$ [29]}),
    .e({\t/a/regfile/regfile$25$ [1],\t/a/regfile/regfile$25$ [29]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1488_o,_al_u1278_o}),
    .q({\t/a/regfile/regfile$25$ [1],\t/a/regfile/regfile$25$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b802|t/a/regfile/reg0_b827  (
    .a({_al_u1256_o,_al_u1319_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .c({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/ID_rs2$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [2],\t/a/regfile/regfile$24$ [27]}),
    .e({\t/a/regfile/regfile$25$ [2],\t/a/regfile/regfile$25$ [27]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1257_o,_al_u1320_o}),
    .q({\t/a/regfile/regfile$25$ [2],\t/a/regfile/regfile$25$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~C*~B*~D*~A+C*~B*~D*~A+C*~B*D*~A+~C*~B*~D*A+C*~B*~D*A+C*~B*D*A"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~C*~B*~D*~A+~C*~B*~D*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b803|t/a/regfile/reg0_b825  (
    .a({open_n39879,_al_u1361_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_16 ,\t/a/ID_rs2$0$_placeOpt_16 }),
    .c({\t/a/ID_rs2$0$_placeOpt_16 ,\t/a/ID_rs2$1$_placeOpt_16 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [3],\t/a/regfile/regfile$24$ [25]}),
    .e({\t/a/regfile/regfile$25$ [3],\t/a/regfile/regfile$25$ [25]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1178_o,_al_u1362_o}),
    .q({\t/a/regfile/regfile$25$ [3],\t/a/regfile/regfile$25$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b804|t/a/regfile/reg0_b824  (
    .a({_al_u1172_o,_al_u1382_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_3 ,\t/a/ID_rs2$0$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$24$ [4],\t/a/ID_rs2$1$_placeOpt_13 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_13 ,\t/a/regfile/regfile$24$ [24]}),
    .e({\t/a/regfile/regfile$25$ [4],\t/a/regfile/regfile$25$ [24]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1173_o,_al_u1383_o}),
    .q({\t/a/regfile/regfile$25$ [4],\t/a/regfile/regfile$25$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b805|t/a/regfile/reg0_b822  (
    .a({_al_u1151_o,_al_u1424_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_2 }),
    .c({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [5],\t/a/regfile/regfile$24$ [22]}),
    .e({\t/a/regfile/regfile$25$ [5],\t/a/regfile/regfile$25$ [22]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1152_o,_al_u1425_o}),
    .q({\t/a/regfile/regfile$25$ [5],\t/a/regfile/regfile$25$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b806|t/a/regfile/reg0_b820  (
    .a({_al_u1130_o,_al_u1466_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_8 ,\t/a/ID_rs2$0$_placeOpt_8 }),
    .c({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [6],\t/a/regfile/regfile$24$ [20]}),
    .e({\t/a/regfile/regfile$25$ [6],\t/a/regfile/regfile$25$ [20]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1131_o,_al_u1467_o}),
    .q({\t/a/regfile/regfile$25$ [6],\t/a/regfile/regfile$25$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~D*~(C*~(0)*~(B)+C*0*~(B)+~(C)*0*B+C*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~D*~(C*~(1)*~(B)+C*1*~(B)+~(C)*1*B+C*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010101000100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b807|t/a/regfile/reg0_b819  (
    .a({_al_u1109_o,_al_u1508_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_16 ,\t/a/ID_rs2$0$_placeOpt_16 }),
    .c({\t/a/regfile/regfile$24$ [7],\t/a/ID_rs2$1$_placeOpt_3 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_3 ,\t/a/regfile/regfile$24$ [19]}),
    .e({\t/a/regfile/regfile$25$ [7],\t/a/regfile/regfile$25$ [19]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1110_o,_al_u1509_o}),
    .q({\t/a/regfile/regfile$25$ [7],\t/a/regfile/regfile$25$ [19]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*~C*D+A*~B*~C*D"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000110011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b808|t/a/regfile/reg0_b818  (
    .a({open_n39955,_al_u1529_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_16 ,\t/a/ID_rs2$0$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$25$ [8],\t/a/ID_rs2$1$_placeOpt_16 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [8],\t/a/regfile/regfile$24$ [18]}),
    .e({\t/a/ID_rs2$0$_placeOpt_1 ,\t/a/regfile/regfile$25$ [18]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1073_o,_al_u1530_o}),
    .q({\t/a/regfile/regfile$25$ [8],\t/a/regfile/regfile$25$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b809|t/a/regfile/reg0_b816  (
    .a({_al_u1067_o,_al_u1571_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .c({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/ID_rs2$1$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [9],\t/a/regfile/regfile$24$ [16]}),
    .e({\t/a/regfile/regfile$25$ [9],\t/a/regfile/regfile$25$ [16]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1068_o,_al_u1572_o}),
    .q({\t/a/regfile/regfile$25$ [9],\t/a/regfile/regfile$25$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+D*~B*C*~A+~D*~B*~C*A+D*~B*~C*A+D*~B*C*A"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("~D*~B*~C*~A+~D*~B*~C*A"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b810|t/a/regfile/reg0_b814  (
    .a({open_n39986,_al_u1613_o}),
    .b({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_8 }),
    .c({\t/a/regfile/regfile$24$ [10],\t/a/ID_rs2$1$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_8 ,\t/a/regfile/regfile$24$ [14]}),
    .e({\t/a/regfile/regfile$25$ [10],\t/a/regfile/regfile$25$ [14]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1682_o,_al_u1614_o}),
    .q({\t/a/regfile/regfile$25$ [10],\t/a/regfile/regfile$25$ [14]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b811|t/a/regfile/reg0_b813  (
    .a({_al_u1676_o,_al_u1634_o}),
    .b({\t/a/ID_rs2$0$_placeOpt_16 ,\t/a/ID_rs2$0$_placeOpt_16 }),
    .c({\t/a/ID_rs2$1$_placeOpt_16 ,\t/a/ID_rs2$1$_placeOpt_16 }),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [11],\t/a/regfile/regfile$24$ [13]}),
    .e({\t/a/regfile/regfile$25$ [11],\t/a/regfile/regfile$25$ [13]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1677_o,_al_u1635_o}),
    .q({\t/a/regfile/regfile$25$ [11],\t/a/regfile/regfile$25$ [13]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b812|t/a/regfile/reg0_b830  (
    .a({\t/a/regfile/regfile$24$ [12],\t/a/ID_rs2$0$_placeOpt_16 }),
    .b({\t/a/ID_rs2$1$_placeOpt_3 ,\t/a/ID_rs2$1$_placeOpt_3 }),
    .c({\t/a/ID_rs2$0$_placeOpt_16 ,\t/a/regfile/regfile$24$ [30]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [12],\t/a/regfile/regfile$25$ [30]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1640_o,_al_u1220_o}),
    .q({\t/a/regfile/regfile$25$ [12],\t/a/regfile/regfile$25$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b815|t/a/regfile/reg0_b828  (
    .a({\t/a/regfile/regfile$24$ [15],\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/regfile/regfile$24$ [28]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [15],\t/a/regfile/regfile$25$ [28]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1577_o,_al_u1283_o}),
    .q({\t/a/regfile/regfile$25$ [15],\t/a/regfile/regfile$25$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b817|t/a/regfile/reg0_b826  (
    .a({\t/a/regfile/regfile$24$ [17],\t/a/ID_rs2$0$_placeOpt_8 }),
    .b({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/ID_rs2$0$_placeOpt_8 ,\t/a/regfile/regfile$24$ [26]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [17],\t/a/regfile/regfile$25$ [26]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1535_o,_al_u1325_o}),
    .q({\t/a/regfile/regfile$25$ [17],\t/a/regfile/regfile$25$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b821|t/a/regfile/reg0_b823  (
    .a({\t/a/regfile/regfile$24$ [21],\t/a/ID_rs2$0$_placeOpt_2 }),
    .b({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/ID_rs2$0$_placeOpt_2 ,\t/a/regfile/regfile$24$ [23]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [21],\t/a/regfile/regfile$25$ [23]}),
    .mi({\t/a/reg_writedat [21],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1430_o,_al_u1388_o}),
    .q({\t/a/regfile/regfile$25$ [21],\t/a/regfile/regfile$25$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*~D*C*~A*B)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*~D*C*~A*B)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000001000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b832|t/a/regfile/reg0_b862  (
    .a({\t/a/WB_rd [0],\t/a/ID_rs1$0$_placeOpt_10 }),
    .b({_al_u256_o,\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$26$ [30]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$27$ [30]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b832_sel_is_3_o ,_al_u519_o}),
    .q({\t/a/regfile/regfile$26$ [0],\t/a/regfile/regfile$26$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~B*~(C*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~B*~(C*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0001001100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0011001100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b833|t/a/regfile/reg0_b860  (
    .a({\t/a/ID_rs1$0$_placeOpt_5 ,\t/a/ID_rs1$0$_placeOpt_5 }),
    .b({\t/a/ID_rs1 [2],\t/a/ID_rs1$1$_placeOpt_5 }),
    .c({\t/a/ID_rs1$1$_placeOpt_5 ,\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [1],\t/a/regfile/regfile$26$ [28]}),
    .e({\t/a/regfile/regfile$27$ [1],\t/a/regfile/regfile$27$ [28]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u771_o,_al_u582_o}),
    .q({\t/a/regfile/regfile$26$ [1],\t/a/regfile/regfile$26$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b834|t/a/regfile/reg0_b858  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1$2$_placeOpt_2 ,\t/a/ID_rs1$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [2],\t/a/regfile/regfile$26$ [26]}),
    .e({\t/a/regfile/regfile$27$ [2],\t/a/regfile/regfile$27$ [26]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u540_o,_al_u624_o}),
    .q({\t/a/regfile/regfile$26$ [2],\t/a/regfile/regfile$26$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~A*~(B*~(C*~(0)*~(D)+C*0*~(D)+~(C)*0*D+C*0*D)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~A*~(B*~(C*~(1)*~(D)+C*1*~(D)+~(C)*1*D+C*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0001000101010001),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0101010101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b835|t/a/regfile/reg0_b857  (
    .a({\t/a/ID_rs1$2$_placeOpt_1 ,\t/a/ID_rs1$0$_placeOpt_2 }),
    .b({\t/a/ID_rs1$1$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$26$ [3],\t/a/ID_rs1$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_2 ,\t/a/regfile/regfile$26$ [25]}),
    .e({\t/a/regfile/regfile$27$ [3],\t/a/regfile/regfile$27$ [25]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u477_o,_al_u645_o}),
    .q({\t/a/regfile/regfile$26$ [3],\t/a/regfile/regfile$26$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b836|t/a/regfile/reg0_b863  (
    .a({\t/a/regfile/regfile$26$ [4],\t/a/ID_rs1$0$_placeOpt_13 }),
    .b({\t/a/regfile/regfile$27$ [4],\t/a/ID_rs1$1$_placeOpt_13 }),
    .c({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/regfile/regfile$26$ [31]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/regfile/regfile$27$ [31]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u442_o,_al_u484_o}),
    .q({\t/a/regfile/regfile$26$ [4],\t/a/regfile/regfile$26$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b837|t/a/regfile/reg0_b856  (
    .a({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/ID_rs1$2$_placeOpt_7 ,\t/a/ID_rs1$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [5],\t/a/regfile/regfile$26$ [24]}),
    .e({\t/a/regfile/regfile$27$ [5],\t/a/regfile/regfile$27$ [24]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u435_o,_al_u666_o}),
    .q({\t/a/regfile/regfile$26$ [5],\t/a/regfile/regfile$26$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b838|t/a/regfile/reg0_b855  (
    .a({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/ID_rs1$2$_placeOpt_7 ,\t/a/ID_rs1$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [6],\t/a/regfile/regfile$26$ [23]}),
    .e({\t/a/regfile/regfile$27$ [6],\t/a/regfile/regfile$27$ [23]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u414_o,_al_u687_o}),
    .q({\t/a/regfile/regfile$26$ [6],\t/a/regfile/regfile$26$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b839|t/a/regfile/reg0_b861  (
    .a({\t/a/regfile/regfile$27$ [7],\t/a/ID_rs1$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$26$ [7],\t/a/ID_rs1$1$_placeOpt_5 }),
    .c({\t/a/ID_rs1$1$_placeOpt_5 ,\t/a/regfile/regfile$26$ [29]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_5 ,\t/a/regfile/regfile$27$ [29]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u379_o,_al_u547_o}),
    .q({\t/a/regfile/regfile$26$ [7],\t/a/regfile/regfile$26$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b840|t/a/regfile/reg0_b853  (
    .a({\t/a/ID_rs1$0$_placeOpt_3 ,\t/a/ID_rs1$0$_placeOpt_3 }),
    .b({\t/a/ID_rs1$1$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$27$ [8],\t/a/ID_rs1$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [8],\t/a/regfile/regfile$26$ [21]}),
    .e({\t/a/ID_rs1$2$_placeOpt_7 ,\t/a/regfile/regfile$27$ [21]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u372_o,_al_u729_o}),
    .q({\t/a/regfile/regfile$26$ [8],\t/a/regfile/regfile$26$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b841|t/a/regfile/reg0_b859  (
    .a({\t/a/regfile/regfile$26$ [9],\t/a/ID_rs1$0$_placeOpt_7 }),
    .b({\t/a/regfile/regfile$27$ [9],\t/a/ID_rs1$1$_placeOpt_7 }),
    .c({\t/a/ID_rs1$1$_placeOpt_7 ,\t/a/regfile/regfile$26$ [27]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_7 ,\t/a/regfile/regfile$27$ [27]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u337_o,_al_u589_o}),
    .q({\t/a/regfile/regfile$26$ [9],\t/a/regfile/regfile$26$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b842|t/a/regfile/reg0_b851  (
    .a({\t/a/ID_rs1$0$_placeOpt_8 ,\t/a/ID_rs1$0$_placeOpt_8 }),
    .b({\t/a/ID_rs1$1$_placeOpt_8 ,\t/a/ID_rs1$1$_placeOpt_8 }),
    .c({\t/a/regfile/regfile$27$ [10],\t/a/ID_rs1$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [10],\t/a/regfile/regfile$26$ [19]}),
    .e({\t/a/ID_rs1$2$_placeOpt_2 ,\t/a/regfile/regfile$27$ [19]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u981_o,_al_u792_o}),
    .q({\t/a/regfile/regfile$26$ [10],\t/a/regfile/regfile$26$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b843|t/a/regfile/reg0_b854  (
    .a({\t/a/regfile/regfile$27$ [11],\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/regfile/regfile$26$ [11],\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/regfile/regfile$26$ [22]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/regfile/regfile$27$ [22]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u946_o,_al_u694_o}),
    .q({\t/a/regfile/regfile$26$ [11],\t/a/regfile/regfile$26$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b844|t/a/regfile/reg0_b849  (
    .a({\t/a/ID_rs1$0$_placeOpt_3 ,\t/a/ID_rs1$0$_placeOpt_3 }),
    .b({\t/a/ID_rs1$1$_placeOpt_3 ,\t/a/ID_rs1$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$27$ [12],\t/a/ID_rs1$2$_placeOpt_7 }),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [12],\t/a/regfile/regfile$26$ [17]}),
    .e({\t/a/ID_rs1$2$_placeOpt_7 ,\t/a/regfile/regfile$27$ [17]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u939_o,_al_u834_o}),
    .q({\t/a/regfile/regfile$26$ [12],\t/a/regfile/regfile$26$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b845|t/a/regfile/reg0_b852  (
    .a({\t/a/regfile/regfile$27$ [13],\t/a/ID_rs1$0$_placeOpt_8 }),
    .b({\t/a/regfile/regfile$26$ [13],\t/a/ID_rs1$1$_placeOpt_8 }),
    .c({\t/a/ID_rs1$1$_placeOpt_8 ,\t/a/regfile/regfile$26$ [20]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_8 ,\t/a/regfile/regfile$27$ [20]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u904_o,_al_u736_o}),
    .q({\t/a/regfile/regfile$26$ [13],\t/a/regfile/regfile$26$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b846|t/a/regfile/reg0_b847  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1$2$_placeOpt_2 ,\t/a/ID_rs1$2$_placeOpt_2 }),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [14],\t/a/regfile/regfile$26$ [15]}),
    .e({\t/a/regfile/regfile$27$ [14],\t/a/regfile/regfile$27$ [15]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u897_o,_al_u876_o}),
    .q({\t/a/regfile/regfile$26$ [14],\t/a/regfile/regfile$26$ [15]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010011000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b848|t/a/regfile/reg0_b850  (
    .a({\t/a/regfile/regfile$26$ [16],\t/a/ID_rs1$0$_placeOpt_8 }),
    .b({\t/a/ID_rs1$1$_placeOpt_8 ,\t/a/ID_rs1$1$_placeOpt_8 }),
    .c({\t/a/ID_rs1$0$_placeOpt_8 ,\t/a/regfile/regfile$26$ [18]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [16],\t/a/regfile/regfile$27$ [18]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u841_o,_al_u799_o}),
    .q({\t/a/regfile/regfile$26$ [16],\t/a/regfile/regfile$26$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*~D*C*B*A)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b864|t/a/regfile/reg0_b895  (
    .a({_al_u256_o,\t/a/ID_rs2$0$_placeOpt_22 }),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2$1$_placeOpt_11 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2$2$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$26$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$27$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b864_sel_is_3_o ,_al_u1214_o}),
    .q({\t/a/regfile/regfile$27$ [0],\t/a/regfile/regfile$27$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~A*~(B*~(C*~(0)*~(D)+C*0*~(D)+~(C)*0*D+C*0*D)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~A*~(B*~(C*~(1)*~(D)+C*1*~(D)+~(C)*1*D+C*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0001000101010001),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0101010101010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b865|t/a/regfile/reg0_b893  (
    .a({\t/a/ID_rs2 [2],\t/a/ID_rs2$0$_placeOpt_4 }),
    .b({\t/a/ID_rs2$1$_placeOpt_1 ,\t/a/ID_rs2$1$_placeOpt_1 }),
    .c({\t/a/regfile/regfile$26$ [1],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/regfile/regfile$26$ [29]}),
    .e({\t/a/regfile/regfile$27$ [1],\t/a/regfile/regfile$27$ [29]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1487_o,_al_u1277_o}),
    .q({\t/a/regfile/regfile$27$ [1],\t/a/regfile/regfile$27$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b866|t/a/regfile/reg0_b891  (
    .a({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/ID_rs2$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [2],\t/a/regfile/regfile$26$ [27]}),
    .e({\t/a/regfile/regfile$27$ [2],\t/a/regfile/regfile$27$ [27]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1256_o,_al_u1319_o}),
    .q({\t/a/regfile/regfile$27$ [2],\t/a/regfile/regfile$27$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*C*~D*~B+A*C*~D*~B+A*C*D*~B+~A*C*~D*B+A*C*~D*B+A*C*D*B"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("~A*C*~D*~B+~A*C*~D*B"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1010000011110000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b867|t/a/regfile/reg0_b878  (
    .a({\t/a/ID_rs2$0$_placeOpt_16 ,\t/a/ID_rs2$0$_placeOpt_16 }),
    .b({open_n40342,\t/a/ID_rs2$1$_placeOpt_16 }),
    .c({\t/a/ID_rs2$1$_placeOpt_16 ,\t/a/ID_rs2$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [3],\t/a/regfile/regfile$26$ [14]}),
    .e({\t/a/regfile/regfile$27$ [3],\t/a/regfile/regfile$27$ [14]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1179_o,_al_u1613_o}),
    .q({\t/a/regfile/regfile$27$ [3],\t/a/regfile/regfile$27$ [14]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b868|t/a/regfile/reg0_b889  (
    .a({\t/a/ID_rs2$0$_placeOpt_3 ,\t/a/ID_rs2$0$_placeOpt_3 }),
    .b({\t/a/ID_rs2$1$_placeOpt_13 ,\t/a/ID_rs2$1$_placeOpt_13 }),
    .c({\t/a/regfile/regfile$27$ [4],\t/a/ID_rs2$2$_placeOpt_6 }),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [4],\t/a/regfile/regfile$26$ [25]}),
    .e({\t/a/ID_rs2$2$_placeOpt_6 ,\t/a/regfile/regfile$27$ [25]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1172_o,_al_u1361_o}),
    .q({\t/a/regfile/regfile$27$ [4],\t/a/regfile/regfile$27$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000011111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b869|t/a/regfile/reg0_b888  (
    .a({\t/a/ID_rs2$0$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_2 }),
    .b({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$26$ [5],\t/a/ID_rs2$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$2$_placeOpt_9 ,\t/a/regfile/regfile$26$ [24]}),
    .e({\t/a/regfile/regfile$27$ [5],\t/a/regfile/regfile$27$ [24]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1151_o,_al_u1382_o}),
    .q({\t/a/regfile/regfile$27$ [5],\t/a/regfile/regfile$27$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~D*~(B*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~D*~(B*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000011111011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b870|t/a/regfile/reg0_b886  (
    .a({\t/a/ID_rs2$0$_placeOpt_2 ,\t/a/ID_rs2$0$_placeOpt_2 }),
    .b({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$26$ [6],\t/a/ID_rs2$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$2$_placeOpt_9 ,\t/a/regfile/regfile$26$ [22]}),
    .e({\t/a/regfile/regfile$27$ [6],\t/a/regfile/regfile$27$ [22]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1130_o,_al_u1424_o}),
    .q({\t/a/regfile/regfile$27$ [6],\t/a/regfile/regfile$27$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b871|t/a/regfile/reg0_b884  (
    .a({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/regfile/regfile$27$ [7],\t/a/ID_rs2$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [7],\t/a/regfile/regfile$26$ [20]}),
    .e({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/regfile/regfile$27$ [20]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1109_o,_al_u1466_o}),
    .q({\t/a/regfile/regfile$27$ [7],\t/a/regfile/regfile$27$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b872|t/a/regfile/reg0_b894  (
    .a({\t/a/regfile/regfile$26$ [8],\t/a/ID_rs2$0$_placeOpt_16 }),
    .b({\t/a/regfile/regfile$27$ [8],\t/a/ID_rs2$1$_placeOpt_3 }),
    .c({\t/a/ID_rs2$0$_placeOpt_16 ,\t/a/regfile/regfile$26$ [30]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_3 ,\t/a/regfile/regfile$27$ [30]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1074_o,_al_u1221_o}),
    .q({\t/a/regfile/regfile$27$ [8],\t/a/regfile/regfile$27$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b873|t/a/regfile/reg0_b883  (
    .a({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/regfile/regfile$27$ [9],\t/a/ID_rs2$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [9],\t/a/regfile/regfile$26$ [19]}),
    .e({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/regfile/regfile$27$ [19]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1067_o,_al_u1508_o}),
    .q({\t/a/regfile/regfile$27$ [9],\t/a/regfile/regfile$27$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0011010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b874|t/a/regfile/reg0_b892  (
    .a({\t/a/regfile/regfile$26$ [10],\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/regfile/regfile$27$ [10],\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/regfile/regfile$26$ [28]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/regfile/regfile$27$ [28]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1683_o,_al_u1284_o}),
    .q({\t/a/regfile/regfile$27$ [10],\t/a/regfile/regfile$27$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b875|t/a/regfile/reg0_b882  (
    .a({\t/a/ID_rs2$0$_placeOpt_1 ,\t/a/ID_rs2$0$_placeOpt_1 }),
    .b({\t/a/ID_rs2$1$_placeOpt_7 ,\t/a/ID_rs2$1$_placeOpt_7 }),
    .c({\t/a/regfile/regfile$27$ [11],\t/a/ID_rs2$2$_placeOpt_8 }),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [11],\t/a/regfile/regfile$26$ [18]}),
    .e({\t/a/ID_rs2$2$_placeOpt_8 ,\t/a/regfile/regfile$27$ [18]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1676_o,_al_u1529_o}),
    .q({\t/a/regfile/regfile$27$ [11],\t/a/regfile/regfile$27$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b876|t/a/regfile/reg0_b890  (
    .a({\t/a/regfile/regfile$27$ [12],\t/a/ID_rs2$0$_placeOpt_8 }),
    .b({\t/a/regfile/regfile$26$ [12],\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/regfile/regfile$26$ [26]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_8 ,\t/a/regfile/regfile$27$ [26]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1641_o,_al_u1326_o}),
    .q({\t/a/regfile/regfile$27$ [12],\t/a/regfile/regfile$27$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*~B*C*~D+A*~B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b1111011110110011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b877|t/a/regfile/reg0_b880  (
    .a({\t/a/ID_rs2$0$_placeOpt_5 ,\t/a/ID_rs2$0$_placeOpt_5 }),
    .b({\t/a/ID_rs2$1$_placeOpt_6 ,\t/a/ID_rs2$1$_placeOpt_6 }),
    .c({\t/a/regfile/regfile$27$ [13],\t/a/ID_rs2$2$_placeOpt_1 }),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [13],\t/a/regfile/regfile$26$ [16]}),
    .e({\t/a/ID_rs2$2$_placeOpt_1 ,\t/a/regfile/regfile$27$ [16]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1634_o,_al_u1571_o}),
    .q({\t/a/regfile/regfile$27$ [13],\t/a/regfile/regfile$27$ [16]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b879|t/a/regfile/reg0_b887  (
    .a({\t/a/regfile/regfile$27$ [15],\t/a/ID_rs2$0$_placeOpt_2 }),
    .b({\t/a/regfile/regfile$26$ [15],\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/regfile/regfile$26$ [23]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_2 ,\t/a/regfile/regfile$27$ [23]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1578_o,_al_u1389_o}),
    .q({\t/a/regfile/regfile$27$ [15],\t/a/regfile/regfile$27$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0001101100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b881|t/a/regfile/reg0_b885  (
    .a({\t/a/ID_rs2$0$_placeOpt_8 ,\t/a/ID_rs2$0$_placeOpt_8 }),
    .b({\t/a/regfile/regfile$26$ [17],\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/regfile/regfile$27$ [17],\t/a/regfile/regfile$26$ [21]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/regfile/regfile$27$ [21]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1536_o,_al_u1431_o}),
    .q({\t/a/regfile/regfile$27$ [17],\t/a/regfile/regfile$27$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b900|t/a/regfile/reg0_b927  (
    .a({\t/a/regfile/regfile$29$ [4],\t/a/ID_rs1$0$_placeOpt_13 }),
    .b({\t/a/regfile/regfile$28$ [4],\t/a/ID_rs1$1$_placeOpt_13 }),
    .c({\t/a/ID_rs1$1$_placeOpt_13 ,\t/a/regfile/regfile$28$ [31]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_13 ,\t/a/regfile/regfile$29$ [31]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u439_o,_al_u481_o}),
    .q({\t/a/regfile/regfile$28$ [4],\t/a/regfile/regfile$28$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b903|t/a/regfile/reg0_b925  (
    .a({\t/a/ID_rs1$0$_placeOpt_19 ,\t/a/ID_rs1$0$_placeOpt_19 }),
    .b({\t/a/regfile/regfile$28$ [7],\t/a/ID_rs1$1$_placeOpt_19 }),
    .c({\t/a/ID_rs1$1$_placeOpt_19 ,\t/a/regfile/regfile$28$ [29]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [7],\t/a/regfile/regfile$29$ [29]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u376_o,_al_u544_o}),
    .q({\t/a/regfile/regfile$28$ [7],\t/a/regfile/regfile$28$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b905|t/a/regfile/reg0_b923  (
    .a({\t/a/regfile/regfile$29$ [9],\t/a/ID_rs1$0$_placeOpt_2 }),
    .b({\t/a/regfile/regfile$28$ [9],\t/a/ID_rs1$1$_placeOpt_2 }),
    .c({\t/a/ID_rs1$1$_placeOpt_2 ,\t/a/regfile/regfile$28$ [27]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_2 ,\t/a/regfile/regfile$29$ [27]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u334_o,_al_u586_o}),
    .q({\t/a/regfile/regfile$28$ [9],\t/a/regfile/regfile$28$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b907|t/a/regfile/reg0_b918  (
    .a({\t/a/regfile/regfile$29$ [11],\t/a/ID_rs1$0$_placeOpt_6 }),
    .b({\t/a/regfile/regfile$28$ [11],\t/a/ID_rs1$1$_placeOpt_6 }),
    .c({\t/a/ID_rs1$1$_placeOpt_6 ,\t/a/regfile/regfile$28$ [22]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_6 ,\t/a/regfile/regfile$29$ [22]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u943_o,_al_u691_o}),
    .q({\t/a/regfile/regfile$28$ [11],\t/a/regfile/regfile$28$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b909|t/a/regfile/reg0_b916  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/regfile/regfile$28$ [13],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [1],\t/a/regfile/regfile$28$ [20]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [13],\t/a/regfile/regfile$29$ [20]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u901_o,_al_u733_o}),
    .q({\t/a/regfile/regfile$28$ [13],\t/a/regfile/regfile$28$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000000110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b912|t/a/regfile/reg0_b914  (
    .a({\t/a/regfile/regfile$28$ [16],\t/a/ID_rs1 [0]}),
    .b({\t/a/regfile/regfile$29$ [16],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [0],\t/a/regfile/regfile$28$ [18]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [1],\t/a/regfile/regfile$29$ [18]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u838_o,_al_u796_o}),
    .q({\t/a/regfile/regfile$28$ [16],\t/a/regfile/regfile$28$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b931|t/a/regfile/reg0_b958  (
    .a({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_4 }),
    .b({\t/a/regfile/regfile$28$ [3],\t/a/ID_rs2$1$_placeOpt_3 }),
    .c({\t/a/ID_rs2$1$_placeOpt_3 ,\t/a/regfile/regfile$28$ [30]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [3],\t/a/regfile/regfile$29$ [30]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1176_o,_al_u1218_o}),
    .q({\t/a/regfile/regfile$29$ [3],\t/a/regfile/regfile$29$ [30]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b936|t/a/regfile/reg0_b956  (
    .a({\t/a/regfile/regfile$28$ [8],\t/a/ID_rs2$0$_placeOpt_16 }),
    .b({\t/a/ID_rs2$1$_placeOpt_3 ,\t/a/ID_rs2$1$_placeOpt_3 }),
    .c({\t/a/ID_rs2$0$_placeOpt_16 ,\t/a/regfile/regfile$28$ [28]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [8],\t/a/regfile/regfile$29$ [28]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1071_o,_al_u1281_o}),
    .q({\t/a/regfile/regfile$29$ [8],\t/a/regfile/regfile$29$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b938|t/a/regfile/reg0_b954  (
    .a({\t/a/regfile/regfile$29$ [10],\t/a/ID_rs2$0$_placeOpt_14 }),
    .b({\t/a/regfile/regfile$28$ [10],\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/regfile/regfile$28$ [26]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_14 ,\t/a/regfile/regfile$29$ [26]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1680_o,_al_u1323_o}),
    .q({\t/a/regfile/regfile$29$ [10],\t/a/regfile/regfile$29$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100001011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b940|t/a/regfile/reg0_b951  (
    .a({\t/a/ID_rs2$0$_placeOpt_18 ,\t/a/ID_rs2$0$_placeOpt_18 }),
    .b({\t/a/regfile/regfile$28$ [12],\t/a/ID_rs2$1$_placeOpt_2 }),
    .c({\t/a/ID_rs2$1$_placeOpt_2 ,\t/a/regfile/regfile$28$ [23]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [12],\t/a/regfile/regfile$29$ [23]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1638_o,_al_u1386_o}),
    .q({\t/a/regfile/regfile$29$ [12],\t/a/regfile/regfile$29$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010100000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b943|t/a/regfile/reg0_b949  (
    .a({\t/a/regfile/regfile$29$ [15],\t/a/ID_rs2$0$_placeOpt_6 }),
    .b({\t/a/regfile/regfile$28$ [15],\t/a/ID_rs2$1$_placeOpt_4 }),
    .c({\t/a/ID_rs2$1$_placeOpt_4 ,\t/a/regfile/regfile$28$ [21]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$0$_placeOpt_6 ,\t/a/regfile/regfile$29$ [21]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1575_o,_al_u1428_o}),
    .q({\t/a/regfile/regfile$29$ [15],\t/a/regfile/regfile$29$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*D*C*~B*A)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b960|t/a/regfile/reg0_b966  (
    .a({_al_u256_o,\t/a/ID_rs1$0$_placeOpt_10 }),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1$1$_placeOpt_10 }),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1$2$_placeOpt_9 }),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$30$ [6]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$31$ [6]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b960_sel_is_3_o ,_al_u412_o}),
    .q({\t/a/regfile/regfile$30$ [0],\t/a/regfile/regfile$30$ [6]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(A*~(B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(A*~(B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0010101000100010),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1010101010100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b961|t/a/regfile/reg0_b965  (
    .a({\t/a/ID_rs1 [2],\t/a/ID_rs1$0$_placeOpt_19 }),
    .b({\t/a/ID_rs1$1$_placeOpt_19 ,\t/a/ID_rs1$1$_placeOpt_19 }),
    .c({\t/a/ID_rs1$0$_placeOpt_19 ,\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [1],\t/a/regfile/regfile$30$ [5]}),
    .e({\t/a/regfile/regfile$31$ [1],\t/a/regfile/regfile$31$ [5]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u769_o,_al_u433_o}),
    .q({\t/a/regfile/regfile$30$ [1],\t/a/regfile/regfile$30$ [5]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(A*~(B*~(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(A*~(B*~(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0010101000100010),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1010101010100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b962|t/a/regfile/reg0_b963  (
    .a({\t/a/ID_rs1 [2],\t/a/ID_rs1$0$_placeOpt_2 }),
    .b({\t/a/ID_rs1$1$_placeOpt_2 ,\t/a/ID_rs1$1$_placeOpt_2 }),
    .c({\t/a/ID_rs1$0$_placeOpt_2 ,\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [2],\t/a/regfile/regfile$30$ [3]}),
    .e({\t/a/regfile/regfile$31$ [2],\t/a/regfile/regfile$31$ [3]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u538_o,_al_u475_o}),
    .q({\t/a/regfile/regfile$30$ [2],\t/a/regfile/regfile$30$ [3]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(A*~(D)*~(C)+A*D*~(C)+~(A)*D*C+A*D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000010011000100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b964|t/a/regfile/reg0_b991  (
    .a({\t/a/regfile/regfile$30$ [4],\t/a/ID_rs1$0$_placeOpt_19 }),
    .b({\t/a/ID_rs1$1$_placeOpt_19 ,\t/a/ID_rs1$1$_placeOpt_19 }),
    .c({\t/a/ID_rs1$0$_placeOpt_19 ,\t/a/regfile/regfile$31$ [31]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$31$ [4],\t/a/regfile/regfile$30$ [31]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u440_o,_al_u482_o}),
    .q({\t/a/regfile/regfile$30$ [4],\t/a/regfile/regfile$30$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0001000010110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b967|t/a/regfile/reg0_b989  (
    .a({\t/a/ID_rs1$0$_placeOpt_19 ,\t/a/ID_rs1$0$_placeOpt_19 }),
    .b({\t/a/regfile/regfile$30$ [7],\t/a/ID_rs1$1$_placeOpt_19 }),
    .c({\t/a/ID_rs1$1$_placeOpt_19 ,\t/a/regfile/regfile$31$ [29]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$31$ [7],\t/a/regfile/regfile$30$ [29]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u377_o,_al_u545_o}),
    .q({\t/a/regfile/regfile$30$ [7],\t/a/regfile/regfile$30$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0010000001110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b969|t/a/regfile/reg0_b987  (
    .a({\t/a/ID_rs1$0$_placeOpt_2 ,\t/a/ID_rs1$0$_placeOpt_2 }),
    .b({\t/a/regfile/regfile$31$ [9],\t/a/ID_rs1$1$_placeOpt_2 }),
    .c({\t/a/ID_rs1$1$_placeOpt_2 ,\t/a/regfile/regfile$31$ [27]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [9],\t/a/regfile/regfile$30$ [27]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u335_o,_al_u587_o}),
    .q({\t/a/regfile/regfile$30$ [9],\t/a/regfile/regfile$30$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0011000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b971|t/a/regfile/reg0_b982  (
    .a({\t/a/regfile/regfile$30$ [11],\t/a/ID_rs1$0$_placeOpt_14 }),
    .b({\t/a/regfile/regfile$31$ [11],\t/a/ID_rs1$1$_placeOpt_14 }),
    .c({\t/a/ID_rs1$1$_placeOpt_14 ,\t/a/regfile/regfile$31$ [22]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1$0$_placeOpt_14 ,\t/a/regfile/regfile$30$ [22]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u944_o,_al_u692_o}),
    .q({\t/a/regfile/regfile$30$ [11],\t/a/regfile/regfile$30$ [22]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b973|t/a/regfile/reg0_b980  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [13],\t/a/regfile/regfile$31$ [20]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [13],\t/a/regfile/regfile$30$ [20]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u902_o,_al_u734_o}),
    .q({\t/a/regfile/regfile$30$ [13],\t/a/regfile/regfile$30$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b976|t/a/regfile/reg0_b978  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [16],\t/a/regfile/regfile$31$ [18]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [16],\t/a/regfile/regfile$30$ [18]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u839_o,_al_u797_o}),
    .q({\t/a/regfile/regfile$30$ [16],\t/a/regfile/regfile$30$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(A*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(A*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000001010000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000011010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b993|t/a/regfile/reg0_b998  (
    .a({\t/a/ID_rs2 [1],\t/a/ID_rs2$0$_placeOpt_10 }),
    .b({\t/a/ID_rs2$0$_placeOpt_10 ,\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2$2$_placeOpt_10 ,\t/a/ID_rs2$2$_placeOpt_10 }),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [1],\t/a/regfile/regfile$30$ [6]}),
    .e({\t/a/regfile/regfile$31$ [1],\t/a/regfile/regfile$31$ [6]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u1485_o,_al_u1128_o}),
    .q({\t/a/regfile/regfile$31$ [1],\t/a/regfile/regfile$31$ [6]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(B*~(D*~(C*~(0)*~(A)+C*0*~(A)+~(C)*0*A+C*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(B*~(D*~(C*~(1)*~(A)+C*1*~(A)+~(C)*1*A+C*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0100000011001100),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1100100011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b994|t/a/regfile/reg0_b997  (
    .a({\t/a/ID_rs2$0$_placeOpt_4 ,\t/a/ID_rs2$0$_placeOpt_4 }),
    .b({\t/a/ID_rs2 [2],\t/a/ID_rs2$1$_placeOpt_3 }),
    .c({\t/a/regfile/regfile$30$ [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2$1$_placeOpt_3 ,\t/a/regfile/regfile$30$ [5]}),
    .e({\t/a/regfile/regfile$31$ [2],\t/a/regfile/regfile$31$ [5]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u1254_o,_al_u1149_o}),
    .q({\t/a/regfile/regfile$31$ [2],\t/a/regfile/regfile$31$ [5]}));  // register.v(63)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_22,control_304}),
    .b({control_23,control_305}),
    .c({\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .f({_al_u3180_o,_al_u3386_o}),
    .q({\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$94$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_reg  (
    .clk(clock_pad),
    .mi({open_n40859,1'b1}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({open_n40865,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r }));  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_reg_placeOpt_1  (
    .clk(clock_pad),
    .mi({open_n40885,1'b1}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({open_n40891,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_1 }));  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_reg_placeOpt_2  (
    .clk(clock_pad),
    .mi({open_n40911,1'b1}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({open_n40917,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_2 }));  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_reg_placeOpt_3  (
    .clk(clock_pad),
    .mi({open_n40937,1'b1}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({open_n40943,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_3 }));  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_reg_placeOpt_4  (
    .clk(clock_pad),
    .mi({open_n40963,1'b1}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({open_n40969,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/dc_r_placeOpt_4 }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({rst_pad,rst_pad}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .q({\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$0$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_25,control_298}),
    .b({control_26,control_299}),
    .c({\trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .f({_al_u3257_o,_al_u3411_o}),
    .q({\trig_node/trigger_node_int_0/U1$1$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_52,control_292}),
    .b({control_53,control_293}),
    .c({\trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u3116_o,_al_u3513_o}),
    .q({\trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$90$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/level_1_r_reg|trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[2],o_data[7]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .q({\trig_node/trigger_node_int_0/U1$10$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_56,control_286}),
    .b({control_55,control_287}),
    .c({\trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .f({_al_u3462_o,_al_u3505_o}),
    .q({\trig_node/trigger_node_int_0/U1$11$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_59,control_280}),
    .b({control_58,control_281}),
    .c({\trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .f({_al_u3133_o,_al_u3266_o}),
    .q({\trig_node/trigger_node_int_0/U1$12$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_62,control_274}),
    .b({control_61,control_275}),
    .c({\trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .f({_al_u3176_o,_al_u3155_o}),
    .q({\trig_node/trigger_node_int_0/U1$13$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_65,control_271}),
    .b({control_64,control_272}),
    .c({\trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .f({_al_u3304_o,_al_u3484_o}),
    .q({\trig_node/trigger_node_int_0/U1$14$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_67,control_262}),
    .b({control_68,control_263}),
    .c({\trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .f({_al_u3450_o,_al_u3270_o}),
    .q({\trig_node/trigger_node_int_0/U1$15$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_71,control_46}),
    .b({control_70,control_47}),
    .c({\trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u3189_o,_al_u3184_o}),
    .q({\trig_node/trigger_node_int_0/U1$16$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_74,control_253}),
    .b({control_73,control_254}),
    .c({\trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .f({_al_u3138_o,_al_u3479_o}),
    .q({\trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[23],o_data[1]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .q({\trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_77,control_244}),
    .b({control_76,control_245}),
    .c({\trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .f({_al_u3291_o,_al_u3142_o}),
    .q({\trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$74$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[22],o_data[22]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .q({\trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$18$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_80,control_43}),
    .b({control_79,control_44}),
    .c({\trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .f({_al_u3441_o,_al_u3428_o}),
    .q({\trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[21],o_data[21]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .q({\trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$19$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_29,control_220}),
    .b({control_28,control_221}),
    .c({\trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .f({_al_u3454_o,_al_u3492_o}),
    .q({\trig_node/trigger_node_int_0/U1$2$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_83,control_214}),
    .b({control_82,control_215}),
    .c({\trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .f({_al_u3300_o,_al_u3244_o}),
    .q({\trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[20],o_data[20]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .q({\trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$20$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_85,control_208}),
    .b({control_86,control_209}),
    .c({\trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .f({_al_u3295_o,_al_u3202_o}),
    .q({\trig_node/trigger_node_int_0/U1$21$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_88,control_178}),
    .b({control_89,control_179}),
    .c({\trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .f({_al_u3172_o,_al_u3437_o}),
    .q({\trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[19],o_data[19]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .q({\trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$22$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_92,control_37}),
    .b({control_91,control_38}),
    .c({\trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u3108_o,_al_u3458_o}),
    .q({\trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[18],o_data[23]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .q({\trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$17$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/level_1_r_reg|trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[18],o_data[5]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .q({\trig_node/trigger_node_int_0/U1$23$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$5$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_94,control_34}),
    .b({control_95,control_35}),
    .c({\trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .f({_al_u3360_o,_al_u3312_o}),
    .q({\trig_node/trigger_node_int_0/U1$24$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101111110011011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_97,control_139}),
    .b({control_98,control_140}),
    .c({\trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .f({_al_u3377_o,_al_u3471_o}),
    .q({\trig_node/trigger_node_int_0/U1$25$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_101,control_31}),
    .b({control_100,control_32}),
    .c({\trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .f({_al_u3364_o,_al_u3308_o}),
    .q({\trig_node/trigger_node_int_0/U1$26$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_103,control_301}),
    .b({control_104,control_302}),
    .c({\trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .f({_al_u3347_o,_al_u3382_o}),
    .q({\trig_node/trigger_node_int_0/U1$27$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTG0(16'b0111011100110011),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/ctl_last_reg  (
    .a({open_n41506,control_106}),
    .b({open_n41507,control_107}),
    .c({open_n41508,\trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({open_n41510,\trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/level_0_r }),
    .e({open_n41511,\trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n41513,\trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .f({open_n41525,_al_u3352_o}),
    .q({open_n41529,\trig_node/trigger_node_int_0/U1$28$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_110,control_289}),
    .b({control_109,control_290}),
    .c({\trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .f({_al_u3373_o,_al_u3394_o}),
    .q({\trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/level_1_r_reg|trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi(o_data[12:11]),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .q({\trig_node/trigger_node_int_0/U1$29$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi(o_data[7:6]),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .q({\trig_node/trigger_node_int_0/U1$3$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$4$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_112,control_283}),
    .b({control_113,control_284}),
    .c({\trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .f({_al_u3223_o,_al_u3509_o}),
    .q({\trig_node/trigger_node_int_0/U1$30$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_115,control_277}),
    .b({control_116,control_278}),
    .c({\trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .f({_al_u3206_o,_al_u3424_o}),
    .q({\trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$85$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[10],o_data[10]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .q({\trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$31$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_118,control_268}),
    .b({control_119,control_269}),
    .c({\trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .f({_al_u3210_o,_al_u3420_o}),
    .q({\trig_node/trigger_node_int_0/U1$32$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_121,control_265}),
    .b({control_122,control_266}),
    .c({\trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .f({_al_u3227_o,_al_u3501_o}),
    .q({\trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[9],i_data[9]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .q({\trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$33$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_125,control_259}),
    .b({control_124,control_260}),
    .c({\trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .f({_al_u3369_o,_al_u3287_o}),
    .q({\trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[8],i_data[8]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .q({\trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$34$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_127,control_256}),
    .b({control_128,control_257}),
    .c({\trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .f({_al_u3253_o,_al_u3496_o}),
    .q({\trig_node/trigger_node_int_0/U1$35$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_130,control_250}),
    .b({control_131,control_251}),
    .c({\trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .f({_al_u3232_o,_al_u3167_o}),
    .q({\trig_node/trigger_node_int_0/U1$36$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_133,control_241}),
    .b({control_134,control_242}),
    .c({\trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .f({_al_u3215_o,_al_u3283_o}),
    .q({\trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[5],i_data[5]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .q({\trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$37$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_136,control_238}),
    .b({control_137,control_239}),
    .c({\trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({_al_u3339_o,_al_u3125_o}),
    .q({\trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[4],i_data[4]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .q({\trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$38$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[3],i_data[3]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .q({\trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$39$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_143,control_235}),
    .b({control_142,control_236}),
    .c({\trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .f({_al_u3475_o,_al_u3121_o}),
    .q({\trig_node/trigger_node_int_0/U1$40$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$71$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_146,control_232}),
    .b({control_145,control_233}),
    .c({\trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({_al_u3343_o,_al_u3399_o}),
    .q({\trig_node/trigger_node_int_0/U1$41$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$70$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_149,control_223}),
    .b({control_148,control_224}),
    .c({\trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .f({_al_u3236_o,_al_u3325_o}),
    .q({\trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[2],i_data[2]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .q({\trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$42$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_151,control_205}),
    .b({control_152,control_206}),
    .c({\trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .f({_al_u3219_o,_al_u3274_o}),
    .q({\trig_node/trigger_node_int_0/U1$43$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$61$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_154,control_202}),
    .b({control_155,control_203}),
    .c({\trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .f({_al_u3317_o,_al_u3488_o}),
    .q({\trig_node/trigger_node_int_0/U1$44$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_157,control_199}),
    .b({control_158,control_200}),
    .c({\trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .f({_al_u3112_o,_al_u3159_o}),
    .q({\trig_node/trigger_node_int_0/U1$45$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$59$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_161,control_196}),
    .b({control_160,control_197}),
    .c({\trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u3193_o,_al_u3416_o}),
    .q({\trig_node/trigger_node_int_0/U1$46$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_163,control_193}),
    .b({control_164,control_194}),
    .c({\trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .f({_al_u3129_o,_al_u3150_o}),
    .q({\trig_node/trigger_node_int_0/U1$47$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$57$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_167,control_190}),
    .b({control_166,control_191}),
    .c({\trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({_al_u3104_o,_al_u3198_o}),
    .q({\trig_node/trigger_node_int_0/U1$48$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$56$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*~(D)*~(C)*~(0)+A*~(B)*~(D)*~(C)*~(0)+A*B*~(D)*~(C)*~(0)+~(A)*~(B)*D*~(C)*~(0)+A*B*D*~(C)*~(0)+~(A)*~(B)*~(D)*C*~(0)+A*~(B)*~(D)*C*~(0)+~(A)*B*~(D)*C*~(0)+A*B*~(D)*C*~(0)+~(A)*~(B)*D*C*~(0)+~(A)*B*D*C*~(0)+A*B*D*C*~(0)+~(A)*~(B)*~(D)*~(C)*0+A*~(B)*~(D)*~(C)*0+~(A)*~(B)*D*~(C)*0+A*~(B)*D*~(C)*0+~(A)*~(B)*~(D)*C*0+A*~(B)*~(D)*C*0+~(A)*B*~(D)*C*0+~(A)*~(B)*D*C*0+A*~(B)*D*C*0+~(A)*B*D*C*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*~(D)*~(C)*~(1)+A*~(B)*~(D)*~(C)*~(1)+A*B*~(D)*~(C)*~(1)+~(A)*~(B)*D*~(C)*~(1)+A*B*D*~(C)*~(1)+~(A)*~(B)*~(D)*C*~(1)+A*~(B)*~(D)*C*~(1)+~(A)*B*~(D)*C*~(1)+A*B*~(D)*C*~(1)+~(A)*~(B)*D*C*~(1)+~(A)*B*D*C*~(1)+A*B*D*C*~(1)+~(A)*~(B)*~(D)*~(C)*1+A*~(B)*~(D)*~(C)*1+~(A)*~(B)*D*~(C)*1+A*~(B)*D*~(C)*1+~(A)*~(B)*~(D)*C*1+A*~(B)*~(D)*C*1+~(A)*B*~(D)*C*1+~(A)*~(B)*D*C*1+A*~(B)*D*C*1+~(A)*B*D*C*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1101100111111011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111001101110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_169,control_187}),
    .b({control_170,control_188}),
    .c({\trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({_al_u3433_o,_al_u3278_o}),
    .q({\trig_node/trigger_node_int_0/U1$49$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_173,control_184}),
    .b({control_172,control_185}),
    .c({\trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({_al_u3467_o,_al_u3146_o}),
    .q({\trig_node/trigger_node_int_0/U1$50$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$54$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("(~(B)*~(A)*~(C)*~(D)*~(0)+B*~(A)*~(C)*~(D)*~(0)+B*A*~(C)*~(D)*~(0)+~(B)*~(A)*C*~(D)*~(0)+B*A*C*~(D)*~(0)+~(B)*~(A)*~(C)*D*~(0)+B*~(A)*~(C)*D*~(0)+~(B)*A*~(C)*D*~(0)+B*A*~(C)*D*~(0)+~(B)*~(A)*C*D*~(0)+~(B)*A*C*D*~(0)+B*A*C*D*~(0)+~(B)*~(A)*~(C)*~(D)*0+B*~(A)*~(C)*~(D)*0+~(B)*~(A)*C*~(D)*0+B*~(A)*C*~(D)*0+~(B)*~(A)*~(C)*D*0+B*~(A)*~(C)*D*0+~(B)*A*~(C)*D*0+~(B)*~(A)*C*D*0+B*~(A)*C*D*0+~(B)*A*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("(~(B)*~(A)*~(C)*~(D)*~(1)+B*~(A)*~(C)*~(D)*~(1)+B*A*~(C)*~(D)*~(1)+~(B)*~(A)*C*~(D)*~(1)+B*A*C*~(D)*~(1)+~(B)*~(A)*~(C)*D*~(1)+B*~(A)*~(C)*D*~(1)+~(B)*A*~(C)*D*~(1)+B*A*~(C)*D*~(1)+~(B)*~(A)*C*D*~(1)+~(B)*A*C*D*~(1)+B*A*C*D*~(1)+~(B)*~(A)*~(C)*~(D)*1+B*~(A)*~(C)*~(D)*1+~(B)*~(A)*C*~(D)*1+B*~(A)*C*~(D)*1+~(B)*~(A)*~(C)*D*1+B*~(A)*~(C)*D*1+~(B)*A*~(C)*D*1+~(B)*~(A)*C*D*1+B*~(A)*C*D*1+~(B)*A*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1011111110011101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b0111011101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/ctl_last_reg|trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/ctl_last_reg  (
    .a({control_176,control_181}),
    .b({control_175,control_182}),
    .c({\trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/ctl_this }),
    .mi({\trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/ctl_this ,\trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 ),
    .f({_al_u3335_o,_al_u3261_o}),
    .q({\trig_node/trigger_node_int_0/U1$51$_ins_detector/ins_detec/ctl_last ,\trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[20],i_data[20]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .q({\trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$52$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[1],i_data[1]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .q({\trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$53$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[18],i_data[18]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .q({\trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$55$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[15],i_data[15]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .q({\trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$58$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[4],o_data[4]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .q({\trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$6$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[13],i_data[13]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .q({\trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$60$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[11],i_data[11]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .q({\trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$62$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[10],i_data[10]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .q({\trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$63$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({i_data[0],i_data[0]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .q({\trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$64$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[9],addr[9]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .q({\trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$65$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[8],addr[8]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .q({\trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$66$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[7],addr[7]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .q({\trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$67$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[6],addr[6]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .q({\trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$68$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[3],o_data[3]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .q({\trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$7$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[31],addr[31]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .q({\trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$72$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[30],addr[30]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .q({\trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$73$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[29],addr[29]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .q({\trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$75$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[28],addr[28]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .q({\trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$76$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[27],addr[27]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .q({\trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$77$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[26],addr[26]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .q({\trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$78$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[25],addr[25]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .q({\trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$79$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[31],o_data[31]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 ),
    .q({\trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$8$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[24],addr[24]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .q({\trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$80$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[23],addr[23]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .q({\trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$81$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[22],addr[22]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .q({\trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$82$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[21],addr[21]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 ),
    .q({\trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$83$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[20],addr[20]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .q({\trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$84$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[19],addr[19]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 ),
    .q({\trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$86$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[18],addr[18]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 ),
    .q({\trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$87$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[17],addr[17]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .q({\trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$88$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[16],addr[16]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 ),
    .q({\trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$89$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({o_data[30],o_data[30]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 ),
    .q({\trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$9$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[14],addr[14]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .q({\trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$91$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[13],addr[13]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .q({\trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$92$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[12],addr[12]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .q({\trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$93$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/level_0_r_reg|trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/level_1_r_reg  (
    .clk(clock_pad),
    .mi({addr[10],addr[10]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 ),
    .q({\trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/level_0_r ,\trig_node/trigger_node_int_0/U1$95$_ins_detector/ins_detec/ctl_this }));  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add0/u0|trig_node/trigger_node_int_0/add0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add0/u0|trig_node/trigger_node_int_0/add0/ucin  (
    .a({\trig_node/trigger_node_int_0/n141 [1],1'b0}),
    .b({1'b1,open_n42962}),
    .f({\trig_node/trigger_node_int_0/force_acq_len [1],open_n42982}),
    .fco(\trig_node/trigger_node_int_0/add0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add0/u0|trig_node/trigger_node_int_0/add0/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add0/u10|trig_node/trigger_node_int_0/add0/u9  (
    .a({\trig_node/trigger_node_int_0/n141 [11],1'b0}),
    .b({1'b0,\trig_node/trigger_node_int_0/n141 [10]}),
    .fci(\trig_node/trigger_node_int_0/add0/c9 ),
    .f(\trig_node/trigger_node_int_0/force_acq_len [11:10]),
    .fco(\trig_node/trigger_node_int_0/add0/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add0/u0|trig_node/trigger_node_int_0/add0/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add0/u12|trig_node/trigger_node_int_0/add0/u11  (
    .a({1'b0,\trig_node/trigger_node_int_0/n141 [12]}),
    .b({\trig_node/trigger_node_int_0/n141 [13],1'b0}),
    .fci(\trig_node/trigger_node_int_0/add0/c11 ),
    .f(\trig_node/trigger_node_int_0/force_acq_len [13:12]),
    .fco(\trig_node/trigger_node_int_0/add0/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add0/u0|trig_node/trigger_node_int_0/add0/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add0/u14|trig_node/trigger_node_int_0/add0/u13  (
    .a(\trig_node/trigger_node_int_0/n141 [15:14]),
    .b(2'b00),
    .fci(\trig_node/trigger_node_int_0/add0/c13 ),
    .f(\trig_node/trigger_node_int_0/force_acq_len [15:14]));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add0/u0|trig_node/trigger_node_int_0/add0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add0/u2|trig_node/trigger_node_int_0/add0/u1  (
    .a(2'b10),
    .b(\trig_node/trigger_node_int_0/n141 [3:2]),
    .fci(\trig_node/trigger_node_int_0/add0/c1 ),
    .f(\trig_node/trigger_node_int_0/force_acq_len [3:2]),
    .fco(\trig_node/trigger_node_int_0/add0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add0/u0|trig_node/trigger_node_int_0/add0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add0/u4|trig_node/trigger_node_int_0/add0/u3  (
    .a({\trig_node/trigger_node_int_0/n141 [5],1'b0}),
    .b({1'b0,\trig_node/trigger_node_int_0/n141 [4]}),
    .fci(\trig_node/trigger_node_int_0/add0/c3 ),
    .f(\trig_node/trigger_node_int_0/force_acq_len [5:4]),
    .fco(\trig_node/trigger_node_int_0/add0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add0/u0|trig_node/trigger_node_int_0/add0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add0/u6|trig_node/trigger_node_int_0/add0/u5  (
    .a({1'b0,\trig_node/trigger_node_int_0/n141 [6]}),
    .b({\trig_node/trigger_node_int_0/n141 [7],1'b0}),
    .fci(\trig_node/trigger_node_int_0/add0/c5 ),
    .f(\trig_node/trigger_node_int_0/force_acq_len [7:6]),
    .fco(\trig_node/trigger_node_int_0/add0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add0/u0|trig_node/trigger_node_int_0/add0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add0/u8|trig_node/trigger_node_int_0/add0/u7  (
    .a(2'b00),
    .b(\trig_node/trigger_node_int_0/n141 [9:8]),
    .fci(\trig_node/trigger_node_int_0/add0/c7 ),
    .f(\trig_node/trigger_node_int_0/force_acq_len [9:8]),
    .fco(\trig_node/trigger_node_int_0/add0/c9 ));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add1/ucin_al_u3549"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add1/u11_al_u3552  (
    .a({\trig_node/trigger_node_int_0/force_acq_reg [13],\trig_node/trigger_node_int_0/force_acq_reg [11]}),
    .b({\trig_node/trigger_node_int_0/force_acq_reg [14],\trig_node/trigger_node_int_0/force_acq_reg [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/add1/c11 ),
    .f({\trig_node/trigger_node_int_0/n179 [13],\trig_node/trigger_node_int_0/n179 [11]}),
    .fco(\trig_node/trigger_node_int_0/add1/c15 ),
    .fx({\trig_node/trigger_node_int_0/n179 [14],\trig_node/trigger_node_int_0/n179 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add1/ucin_al_u3549"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add1/u15_al_u3553  (
    .a({open_n43160,\trig_node/trigger_node_int_0/force_acq_reg [15]}),
    .c(2'b00),
    .d({open_n43165,1'b0}),
    .fci(\trig_node/trigger_node_int_0/add1/c15 ),
    .f({open_n43182,\trig_node/trigger_node_int_0/n179 [15]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add1/ucin_al_u3549"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add1/u3_al_u3550  (
    .a({\trig_node/trigger_node_int_0/force_acq_reg [5],\trig_node/trigger_node_int_0/force_acq_reg [3]}),
    .b({\trig_node/trigger_node_int_0/force_acq_reg [6],\trig_node/trigger_node_int_0/force_acq_reg [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/add1/c3 ),
    .f({\trig_node/trigger_node_int_0/n179 [5],\trig_node/trigger_node_int_0/n179 [3]}),
    .fco(\trig_node/trigger_node_int_0/add1/c7 ),
    .fx({\trig_node/trigger_node_int_0/n179 [6],\trig_node/trigger_node_int_0/n179 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add1/ucin_al_u3549"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/add1/u7_al_u3551  (
    .a({\trig_node/trigger_node_int_0/force_acq_reg [9],\trig_node/trigger_node_int_0/force_acq_reg [7]}),
    .b({\trig_node/trigger_node_int_0/force_acq_reg [10],\trig_node/trigger_node_int_0/force_acq_reg [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/add1/c7 ),
    .f({\trig_node/trigger_node_int_0/n179 [9],\trig_node/trigger_node_int_0/n179 [7]}),
    .fco(\trig_node/trigger_node_int_0/add1/c11 ),
    .fx({\trig_node/trigger_node_int_0/n179 [10],\trig_node/trigger_node_int_0/n179 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/add1/ucin_al_u3549"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/add1/ucin_al_u3549  (
    .a({\trig_node/trigger_node_int_0/force_acq_reg [1],1'b0}),
    .b({\trig_node/trigger_node_int_0/force_acq_reg [2],\trig_node/trigger_node_int_0/force_acq_reg [0]}),
    .c(2'b00),
    .ce(\trig_node/trigger_node_int_0/n177 ),
    .clk(clock_pad),
    .d(2'b01),
    .e(2'b01),
    .mi(\trig_node/trigger_node_int_0/n179 [1:0]),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .f({\trig_node/trigger_node_int_0/n179 [1],open_n43236}),
    .fco(\trig_node/trigger_node_int_0/add1/c3 ),
    .fx({\trig_node/trigger_node_int_0/n179 [2],\trig_node/trigger_node_int_0/n179 [0]}),
    .q(\trig_node/trigger_node_int_0/force_acq_reg [1:0]));
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~A*~D*~C*~B+A*~D*~C*~B+~A*D*~C*~B+A*D*~C*~B+~A*~D*C*~B+A*~D*C*~B+~A*D*C*~B+A*D*C*~B+~A*~D*~C*B+A*~D*~C*B+~A*D*~C*B+A*D*~C*B+~A*~D*C*B+A*~D*C*B+~A*D*C*B+A*D*C*B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0011001100110011),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/force_acq_fin_reg|trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last_reg  (
    .a({open_n43237,control_310}),
    .b({\trig_node/trigger_node_int_0/n177 ,control_311}),
    .c({open_n43238,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({open_n43240,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n43242,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .f({open_n43254,_al_u3390_o}),
    .q({\trig_node/trigger_node_int_0/force_acq_fin ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last }));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/force_acq_fin_reg|trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last_reg_placeOpt_1  (
    .a({open_n43258,control_310}),
    .b({open_n43259,control_311}),
    .c({\trig_node/trigger_node_int_0/n177 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({open_n43261,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/force_acq_fin ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n43263,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,open_n43280}));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*~D+A*B*C*~D+A*~B*~C*D+A*B*~C*D+A*~B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1111111111111111),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1010101010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/force_acq_fin_reg|trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last_reg_placeOpt_2  (
    .a({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,control_310}),
    .b({open_n43281,control_311}),
    .c({open_n43282,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({open_n43284,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/n177 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n43286,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_2 ,open_n43303}));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1100111111001111),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1100111111001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/force_acq_fin_reg|trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last_reg_placeOpt_3  (
    .a({open_n43304,control_310}),
    .b({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,control_311}),
    .c({\trig_node/trigger_node_int_0/n177 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({open_n43306,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r }),
    .e({open_n43307,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n43309,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_3 ,open_n43326}));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1111010111110101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1111010111110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/force_acq_fin_reg|trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last_reg_placeOpt_4  (
    .a({\trig_node/trigger_node_int_0/n177 ,control_310}),
    .b({open_n43327,control_311}),
    .c({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({open_n43329,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r }),
    .e({open_n43330,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n43332,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_4 ,open_n43349}));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0000111100001111),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/force_acq_fin_reg|trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last_reg_placeOpt_5  (
    .a({open_n43350,control_310}),
    .b({open_n43351,control_311}),
    .c({\trig_node/trigger_node_int_0/n177 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({open_n43353,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n43355,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_5 ,open_n43372}));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~D*~B*~C*~A+D*~B*~C*~A+~D*B*~C*~A+D*B*~C*~A+~D*~B*C*~A+D*~B*C*~A+~D*B*C*~A+D*B*C*~A+~D*~B*~C*A+D*~B*~C*A+~D*B*~C*A+D*B*~C*A+~D*~B*C*A+D*~B*C*A+~D*B*C*A+D*B*C*A"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0101010101010101),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/force_acq_fin_reg|trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last_reg_placeOpt_6  (
    .a({\trig_node/trigger_node_int_0/n177 ,control_310}),
    .b({open_n43373,control_311}),
    .c({open_n43374,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({open_n43376,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n43378,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_6 ,open_n43395}));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*~C*D+A*~B*~C*D+~A*B*~C*D+A*B*~C*D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~A*B*~C*~D+A*B*~C*~D+~A*B*C*~D+A*B*C*~D+~A*B*~C*D+A*B*~C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1111111111111111),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1100110011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/force_acq_fin_reg|trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last_reg_placeOpt_7  (
    .a({open_n43396,control_310}),
    .b({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,control_311}),
    .c({open_n43397,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({open_n43399,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/n177 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n43401,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_7 ,open_n43418}));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~A*~B*~C*~D+A*~B*~C*~D+~A*B*~C*~D+A*B*~C*~D+~A*~B*C*~D+A*~B*C*~D+~A*B*C*~D+A*B*C*~D+~A*~B*C*D+A*~B*C*D+~A*B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b1111000011111111),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1111000011111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/force_acq_fin_reg|trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last_reg_placeOpt_8  (
    .a({open_n43419,control_310}),
    .b({open_n43420,control_311}),
    .c({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/n177 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r }),
    .e({open_n43422,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n43424,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_8 ,open_n43441}));  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\detecEdge.v(41)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*~(C)*~(D)*~(0)+A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+~(A)*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*D*~(0)+A*~(B)*~(C)*D*~(0)+~(A)*B*~(C)*D*~(0)+A*B*~(C)*D*~(0)+~(A)*~(B)*C*D*~(0)+~(A)*B*C*D*~(0)+A*B*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+A*~(B)*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*B*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0+~(A)*B*C*D*0)"),
    //.LUTF1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C"),
    //.LUTG0("(~(A)*~(B)*~(C)*~(D)*~(1)+A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+~(A)*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*D*~(1)+A*~(B)*~(C)*D*~(1)+~(A)*B*~(C)*D*~(1)+A*B*~(C)*D*~(1)+~(A)*~(B)*C*D*~(1)+~(A)*B*C*D*~(1)+A*B*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+A*~(B)*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*B*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1+~(A)*B*C*D*1)"),
    //.LUTG1("~A*~B*~D*~C+A*~B*~D*~C+~A*B*~D*~C+A*B*~D*~C+~A*~B*D*~C+A*~B*D*~C+~A*B*D*~C+A*B*D*~C+~A*~B*~D*C+A*~B*~D*C+~A*B*~D*C+A*B*~D*C+~A*~B*D*C+A*~B*D*C+~A*B*D*C+A*B*D*C"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101111110011011),
    .INIT_LUTF1(16'b0000000011111111),
    .INIT_LUTG0(16'b0111011100110011),
    .INIT_LUTG1(16'b1111111111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/force_acq_fin_reg|trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last_reg_placeOpt_9  (
    .a({open_n43442,control_310}),
    .b({open_n43443,control_311}),
    .c({open_n43444,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_last }),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/n177 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/level_0_r }),
    .e({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_1 ,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .mi({open_n43447,\trig_node/trigger_node_int_0/U1$96$_ins_detector/ins_detec/ctl_this }),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync ),
    .q({\trig_node/trigger_node_int_0/force_acq_fin_placeOpt_9 ,open_n43464}));  // D:/td/td/cw\detecEdge.v(41)
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/ucin_al_u3554"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/u11_al_u3557  (
    .a({status_13,status_11}),
    .b({status_14,status_12}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c11 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [13],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [11]}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c15 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [14],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/ucin_al_u3554"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/u15_al_u3558  (
    .a({open_n43483,status_15}),
    .c(2'b00),
    .d({open_n43488,1'b0}),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c15 ),
    .f({open_n43505,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [15]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/ucin_al_u3554"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/u3_al_u3555  (
    .a({status_5,status_3}),
    .b({status_6,status_4}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c3 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [5],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [3]}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c7 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [6],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/ucin_al_u3554"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/u7_al_u3556  (
    .a({status_9,status_7}),
    .b({status_10,status_8}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c7 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [9],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [7]}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c11 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [10],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/ucin_al_u3554"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/ucin_al_u3554  (
    .a({status_1,1'b0}),
    .b({status_2,status_0}),
    .c(2'b00),
    .clk(clock_pad),
    .d(2'b01),
    .e(2'b01),
    .mi({status_1,status_0}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [1],open_n43560}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add0/c3 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [2],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [0]}),
    .q(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [1:0]));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/ucin_al_u3559"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/u11_al_u3562  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [13],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [11]}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [14],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c11 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [13],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [11]}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c15 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [14],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/ucin_al_u3559"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/u15_al_u3563  (
    .a({open_n43579,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [15]}),
    .c(2'b00),
    .d({open_n43584,1'b0}),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c15 ),
    .f({open_n43601,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [15]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/ucin_al_u3559"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/u3_al_u3560  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [5],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [3]}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [6],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c3 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [5],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [3]}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c7 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [6],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/ucin_al_u3559"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/u7_al_u3561  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [9],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [7]}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [10],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c7 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [9],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [7]}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c11 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [10],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/ucin_al_u3559"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/ucin_al_u3559  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [1],1'b0}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [2],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [0]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [1],open_n43660}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/add1/c3 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [2],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_cin  (
    .a(2'b01),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [0],open_n43663}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_10|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_9  (
    .a(2'b00),
    .b(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [10:9]),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c9 ),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_12|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_11  (
    .a(2'b00),
    .b(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [12:11]),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c11 ),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_14|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_13  (
    .a(2'b00),
    .b(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [14:13]),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c13 ),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_2|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_1  (
    .a(2'b01),
    .b(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [2:1]),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c1 ),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_4|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_3  (
    .a(2'b01),
    .b(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [4:3]),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c3 ),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_6|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_5  (
    .a(2'b01),
    .b(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [6:5]),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c5 ),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_8|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_7  (
    .a(2'b00),
    .b(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [8:7]),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c7 ),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_cout|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_15  (
    .a(2'b00),
    .b({1'b1,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [15]}),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/lt0_c15 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n19 ,open_n43875}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/overflow_reg  (
    .a({_al_u3081_o,_al_u3081_o}),
    .b({_al_u3083_o,_al_u3083_o}),
    .c({_al_u3085_o,_al_u3085_o}),
    .clk(clock_pad),
    .d({_al_u3086_o,_al_u3086_o}),
    .mi({open_n43892,status_16}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({open_n43898,status_16}));  // D:/td/td/cw\write_ctrl.v(50)
  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~C)*~(~0*B))"),
    //.LUTF1("~A*~B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*~B*~C*D+A*~B*C*D+A*B*C*D"),
    //.LUTG0("(A*~(D*~C)*~(~1*B))"),
    //.LUTG1("~A*~B*~C*~D+~A*~B*C*~D+~A*B*C*~D+A*~B*~C*D+A*~B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000100010),
    .INIT_LUTF1(16'b1010001001010001),
    .INIT_LUTG0(16'b1010000010101010),
    .INIT_LUTG1(16'b1010001001010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b14|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b12  (
    .a({status_3,_al_u3055_o}),
    .b({status_14,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [14]}),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [14],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [12]}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [3],status_12}),
    .e({open_n43900,status_14}),
    .mi({status_14,status_12}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3065_o,_al_u3056_o}),
    .q({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [14],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [12]}));  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\write_ctrl.v(42)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("~A*~B*~C*~D+~A*B*~C*~D+~A*~B*C*D+~A*B*C*D"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("A*~B*~C*~D+A*B*~C*~D+A*~B*C*D+A*B*C*D"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0101000000000101),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1010000000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b3|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg0_b5  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [3],_al_u3064_o}),
    .b({open_n43916,_al_u3065_o}),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [5],_al_u3066_o}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [5],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [5]}),
    .e({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [3],status_5}),
    .mi({status_3,status_5}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .f({_al_u3075_o,_al_u3067_o}),
    .q({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [3],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/addr_tmp [5]}));  // D:/td/td/cw\write_ctrl.v(42)
  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    //.LUT1("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010111000),
    .INIT_LUT1(16'b0000000010111000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b9  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [0],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [9]}),
    .b({\trig_node/trigger_node_int_0/emb_store_en ,\trig_node/trigger_node_int_0/emb_store_en }),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [0],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [9]}),
    .clk(clock_pad),
    .d({status_17,status_17}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [0],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [9]}));  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    //.LUT1("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010111000),
    .INIT_LUT1(16'b0000000010111000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b10|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b8  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [10],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [8]}),
    .b({\trig_node/trigger_node_int_0/emb_store_en ,\trig_node/trigger_node_int_0/emb_store_en }),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [10],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [8]}),
    .clk(clock_pad),
    .d({status_17,status_17}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [10],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [8]}));  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    //.LUT1("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010111000),
    .INIT_LUT1(16'b0000000010111000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b11|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b7  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [11],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [7]}),
    .b({\trig_node/trigger_node_int_0/emb_store_en ,\trig_node/trigger_node_int_0/emb_store_en }),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [11],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [7]}),
    .clk(clock_pad),
    .d({status_17,status_17}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [11],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [7]}));  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    //.LUT1("(~D*(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010111000),
    .INIT_LUT1(16'b0000000011011000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b12|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b6  (
    .a({\trig_node/trigger_node_int_0/emb_store_en ,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [6]}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [12],\trig_node/trigger_node_int_0/emb_store_en }),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [12],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [6]}),
    .clk(clock_pad),
    .d({status_17,status_17}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [12],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [6]}));  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    //.LUT1("(~C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010111000),
    .INIT_LUT1(16'b0000110100001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b13|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b5  (
    .a({\trig_node/trigger_node_int_0/emb_store_en ,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [5]}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [13],\trig_node/trigger_node_int_0/emb_store_en }),
    .c({status_17,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [5]}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [13],status_17}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [13],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [5]}));  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    //.LUT1("(~C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010111000),
    .INIT_LUT1(16'b0000101100001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b14|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b4  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [14],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [4]}),
    .b({\trig_node/trigger_node_int_0/emb_store_en ,\trig_node/trigger_node_int_0/emb_store_en }),
    .c({status_17,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [4]}),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [14],status_17}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [14],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [4]}));  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    //.LUT1("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010111000),
    .INIT_LUT1(16'b0000000010111000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b15|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b3  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [15],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [3]}),
    .b({\trig_node/trigger_node_int_0/emb_store_en ,\trig_node/trigger_node_int_0/emb_store_en }),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [15],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [3]}),
    .clk(clock_pad),
    .d({status_17,status_17}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [15],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [3]}));  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(67)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B))"),
    //.LUT1("(~D*(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010111000),
    .INIT_LUT1(16'b0000000011011000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b1|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg1_b2  (
    .a({\trig_node/trigger_node_int_0/emb_store_en ,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [2]}),
    .b({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n16 [1],\trig_node/trigger_node_int_0/emb_store_en }),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [1],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [2]}),
    .clk(clock_pad),
    .d({status_17,status_17}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [1],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/stop_count [2]}));  // D:/td/td/cw\write_ctrl.v(67)
  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~B)"),
    //.LUT1("(D*~B)"),
    .CEMUX("CE"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001000100010),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b0|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b2  (
    .a({open_n44077,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [2]}),
    .b({_al_u3069_o,_al_u3069_o}),
    .ce(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13$0$_en ),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [0],open_n44080}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({status_0,status_2}));  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~B)"),
    //.LUT1("(D*~B)"),
    .CEMUX("CE"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001000100010),
    .INIT_LUT1(16'b0011001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b10|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b5  (
    .a({open_n44098,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [5]}),
    .b({_al_u3069_o,_al_u3069_o}),
    .ce(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13$0$_en ),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [10],open_n44101}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({status_10,status_5}));  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~A)"),
    //.LUT1("(D*~A)"),
    .CEMUX("CE"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010100000000),
    .INIT_LUT1(16'b0101010100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b11|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b4  (
    .a({_al_u3069_o,_al_u3069_o}),
    .ce(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13$0$_en ),
    .clk(clock_pad),
    .d({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [11],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [4]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({status_11,status_4}));  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~B)"),
    //.LUT1("(A*~B)"),
    .CEMUX("CE"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001000100010),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b12|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b3  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [12],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [3]}),
    .b({_al_u3069_o,_al_u3069_o}),
    .ce(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13$0$_en ),
    .clk(clock_pad),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({status_12,status_3}));  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~B)"),
    //.LUT1("(C*~B)"),
    .CEMUX("CE"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010001000100010),
    .INIT_LUT1(16'b0011000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b13|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b1  (
    .a({open_n44161,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [1]}),
    .b({_al_u3069_o,_al_u3069_o}),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [13],open_n44162}),
    .ce(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13$0$_en ),
    .clk(clock_pad),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({status_13,status_1}));  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~A)"),
    //.LUT1("(C*~A)"),
    .CEMUX("CE"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010100000000),
    .INIT_LUT1(16'b0101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b14|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b9  (
    .a({_al_u3069_o,_al_u3069_o}),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [14],open_n44184}),
    .ce(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13$0$_en ),
    .clk(clock_pad),
    .d({open_n44185,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [9]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({status_14,status_9}));  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~B)"),
    //.LUT1("(A*~B)"),
    .CEMUX("CE"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011001100000000),
    .INIT_LUT1(16'b0010001000100010),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b15|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b8  (
    .a({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [15],open_n44203}),
    .b({_al_u3069_o,_al_u3069_o}),
    .ce(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13$0$_en ),
    .clk(clock_pad),
    .d({open_n44206,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [8]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({status_15,status_8}));  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  // D:/td/td/cw\write_ctrl.v(59)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("INV"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011001100),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b6|trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/reg2_b7  (
    .b({open_n44226,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [7]}),
    .c({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13 [6],open_n44227}),
    .ce(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n13$0$_en ),
    .clk(clock_pad),
    .d({_al_u3069_o,_al_u3069_o}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 ),
    .q({status_6,status_7}));  // D:/td/td/cw\write_ctrl.v(59)
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/ucin_al_u3564"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/u11_al_u3567  (
    .a({control_19,control_17}),
    .b({control_20,control_18}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c11 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [13],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [11]}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c15 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [14],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/ucin_al_u3564"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/u15_al_u3568  (
    .a({open_n44263,control_21}),
    .c(2'b11),
    .d({open_n44268,1'b0}),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c15 ),
    .f({open_n44285,\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [15]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/ucin_al_u3564"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/u3_al_u3565  (
    .a({control_11,control_9}),
    .b({control_12,control_10}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c3 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [5],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [3]}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c7 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [6],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/ucin_al_u3564"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/u7_al_u3566  (
    .a({control_15,control_13}),
    .b({control_16,control_14}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c7 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [9],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [7]}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c11 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [10],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/ucin_al_u3564"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/ucin_al_u3564  (
    .a({control_7,1'b0}),
    .b({control_8,control_6}),
    .c(2'b11),
    .ce(jupdate),
    .clk(jtck),
    .d(2'b01),
    .e(2'b01),
    .mi(\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [8:7]),
    .sr(\cfg_int/wrapper_cfg_inst/rst_placeOpt_15 ),
    .f({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [1],open_n44339}),
    .fco(\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/sub0/c3 ),
    .fx({\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [2],\trig_node/trigger_node_int_0/ins_emb_ctrl/ins_wt_ctrl/n4 [0]}),
    .q({control_8,control_7}));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/lt0_0|trig_node/trigger_node_int_0/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/lt0_0|trig_node/trigger_node_int_0/lt0_cin  (
    .a({\trig_node/trigger_node_int_0/force_acq_reg [0],1'b0}),
    .b({\trig_node/trigger_node_int_0/force_acq_len [0],open_n44340}),
    .fco(\trig_node/trigger_node_int_0/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/lt0_0|trig_node/trigger_node_int_0/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/lt0_10|trig_node/trigger_node_int_0/lt0_9  (
    .a(\trig_node/trigger_node_int_0/force_acq_reg [10:9]),
    .b(\trig_node/trigger_node_int_0/force_acq_len [10:9]),
    .fci(\trig_node/trigger_node_int_0/lt0_c9 ),
    .fco(\trig_node/trigger_node_int_0/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/lt0_0|trig_node/trigger_node_int_0/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/lt0_12|trig_node/trigger_node_int_0/lt0_11  (
    .a(\trig_node/trigger_node_int_0/force_acq_reg [12:11]),
    .b(\trig_node/trigger_node_int_0/force_acq_len [12:11]),
    .fci(\trig_node/trigger_node_int_0/lt0_c11 ),
    .fco(\trig_node/trigger_node_int_0/lt0_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/lt0_0|trig_node/trigger_node_int_0/lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/lt0_14|trig_node/trigger_node_int_0/lt0_13  (
    .a(\trig_node/trigger_node_int_0/force_acq_reg [14:13]),
    .b(\trig_node/trigger_node_int_0/force_acq_len [14:13]),
    .fci(\trig_node/trigger_node_int_0/lt0_c13 ),
    .fco(\trig_node/trigger_node_int_0/lt0_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/lt0_0|trig_node/trigger_node_int_0/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/lt0_2|trig_node/trigger_node_int_0/lt0_1  (
    .a(\trig_node/trigger_node_int_0/force_acq_reg [2:1]),
    .b(\trig_node/trigger_node_int_0/force_acq_len [2:1]),
    .fci(\trig_node/trigger_node_int_0/lt0_c1 ),
    .fco(\trig_node/trigger_node_int_0/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/lt0_0|trig_node/trigger_node_int_0/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/lt0_4|trig_node/trigger_node_int_0/lt0_3  (
    .a(\trig_node/trigger_node_int_0/force_acq_reg [4:3]),
    .b(\trig_node/trigger_node_int_0/force_acq_len [4:3]),
    .fci(\trig_node/trigger_node_int_0/lt0_c3 ),
    .fco(\trig_node/trigger_node_int_0/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/lt0_0|trig_node/trigger_node_int_0/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/lt0_6|trig_node/trigger_node_int_0/lt0_5  (
    .a(\trig_node/trigger_node_int_0/force_acq_reg [6:5]),
    .b(\trig_node/trigger_node_int_0/force_acq_len [6:5]),
    .fci(\trig_node/trigger_node_int_0/lt0_c5 ),
    .fco(\trig_node/trigger_node_int_0/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/lt0_0|trig_node/trigger_node_int_0/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/lt0_8|trig_node/trigger_node_int_0/lt0_7  (
    .a(\trig_node/trigger_node_int_0/force_acq_reg [8:7]),
    .b(\trig_node/trigger_node_int_0/force_acq_len [8:7]),
    .fci(\trig_node/trigger_node_int_0/lt0_c7 ),
    .fco(\trig_node/trigger_node_int_0/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/lt0_0|trig_node/trigger_node_int_0/lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/lt0_cout|trig_node/trigger_node_int_0/lt0_15  (
    .a({1'b0,\trig_node/trigger_node_int_0/force_acq_reg [15]}),
    .b({1'b1,\trig_node/trigger_node_int_0/force_acq_len [15]}),
    .fci(\trig_node/trigger_node_int_0/lt0_c15 ),
    .f({\trig_node/trigger_node_int_0/n177 ,open_n44552}));
  // D:/td/td/cw\trigger_node.v(87)
  // D:/td/td/cw\trigger_node.v(86)
  EG_PHY_MSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/pause_sync0_reg|trig_node/trigger_node_int_0/pause_sync_reg  (
    .clk(clock_pad),
    .mi({control_1,\trig_node/trigger_node_int_0/pause_sync0 }),
    .q({\trig_node/trigger_node_int_0/pause_sync0 ,\trig_node/trigger_node_int_0/pause_sync }));  // D:/td/td/cw\trigger_node.v(87)
  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/reg0_b10|trig_node/trigger_node_int_0/reg0_b9  (
    .ce(\trig_node/trigger_node_int_0/n177 ),
    .clk(clock_pad),
    .mi(\trig_node/trigger_node_int_0/n179 [10:9]),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .q(\trig_node/trigger_node_int_0/force_acq_reg [10:9]));  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/reg0_b11|trig_node/trigger_node_int_0/reg0_b8  (
    .ce(\trig_node/trigger_node_int_0/n177 ),
    .clk(clock_pad),
    .mi({\trig_node/trigger_node_int_0/n179 [11],\trig_node/trigger_node_int_0/n179 [8]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .q({\trig_node/trigger_node_int_0/force_acq_reg [11],\trig_node/trigger_node_int_0/force_acq_reg [8]}));  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/reg0_b12|trig_node/trigger_node_int_0/reg0_b7  (
    .ce(\trig_node/trigger_node_int_0/n177 ),
    .clk(clock_pad),
    .mi({\trig_node/trigger_node_int_0/n179 [12],\trig_node/trigger_node_int_0/n179 [7]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .q({\trig_node/trigger_node_int_0/force_acq_reg [12],\trig_node/trigger_node_int_0/force_acq_reg [7]}));  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/reg0_b13|trig_node/trigger_node_int_0/reg0_b6  (
    .ce(\trig_node/trigger_node_int_0/n177 ),
    .clk(clock_pad),
    .mi({\trig_node/trigger_node_int_0/n179 [13],\trig_node/trigger_node_int_0/n179 [6]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .q({\trig_node/trigger_node_int_0/force_acq_reg [13],\trig_node/trigger_node_int_0/force_acq_reg [6]}));  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/reg0_b14|trig_node/trigger_node_int_0/reg0_b5  (
    .ce(\trig_node/trigger_node_int_0/n177 ),
    .clk(clock_pad),
    .mi({\trig_node/trigger_node_int_0/n179 [14],\trig_node/trigger_node_int_0/n179 [5]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .q({\trig_node/trigger_node_int_0/force_acq_reg [14],\trig_node/trigger_node_int_0/force_acq_reg [5]}));  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/reg0_b15|trig_node/trigger_node_int_0/reg0_b4  (
    .ce(\trig_node/trigger_node_int_0/n177 ),
    .clk(clock_pad),
    .mi({\trig_node/trigger_node_int_0/n179 [15],\trig_node/trigger_node_int_0/n179 [4]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .q({\trig_node/trigger_node_int_0/force_acq_reg [15],\trig_node/trigger_node_int_0/force_acq_reg [4]}));  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_MSLICE #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \trig_node/trigger_node_int_0/reg0_b2|trig_node/trigger_node_int_0/reg0_b3  (
    .ce(\trig_node/trigger_node_int_0/n177 ),
    .clk(clock_pad),
    .mi({\trig_node/trigger_node_int_0/n179 [2],\trig_node/trigger_node_int_0/n179 [3]}),
    .sr(\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 ),
    .q({\trig_node/trigger_node_int_0/force_acq_reg [2],\trig_node/trigger_node_int_0/force_acq_reg [3]}));  // D:/td/td/cw\trigger_node.v(122)
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/sub0/u0|trig_node/trigger_node_int_0/sub0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("SR"))
    \trig_node/trigger_node_int_0/sub0/u0|trig_node/trigger_node_int_0/sub0/ucin  (
    .a({control_6,1'b0}),
    .b({1'b0,open_n44744}),
    .ce(jupdate),
    .clk(jtck),
    .mi({open_n44759,\cfg_int/wrapper_cfg_inst/reg_inst/cshift_r [6]}),
    .sr(\cfg_int/wrapper_cfg_inst/rst ),
    .f({\trig_node/trigger_node_int_0/force_acq_len [0],open_n44760}),
    .fco(\trig_node/trigger_node_int_0/sub0/c1 ),
    .q({open_n44763,control_6}));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/sub0/u0|trig_node/trigger_node_int_0/sub0/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/sub0/u10|trig_node/trigger_node_int_0/sub0/u9  (
    .a({control_16,control_15}),
    .b(2'b00),
    .fci(\trig_node/trigger_node_int_0/sub0/c9 ),
    .f(\trig_node/trigger_node_int_0/n141 [10:9]),
    .fco(\trig_node/trigger_node_int_0/sub0/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/sub0/u0|trig_node/trigger_node_int_0/sub0/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/sub0/u12|trig_node/trigger_node_int_0/sub0/u11  (
    .a({control_18,control_17}),
    .b(2'b00),
    .fci(\trig_node/trigger_node_int_0/sub0/c11 ),
    .f(\trig_node/trigger_node_int_0/n141 [12:11]),
    .fco(\trig_node/trigger_node_int_0/sub0/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/sub0/u0|trig_node/trigger_node_int_0/sub0/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/sub0/u14|trig_node/trigger_node_int_0/sub0/u13  (
    .a({control_20,control_19}),
    .b(2'b00),
    .fci(\trig_node/trigger_node_int_0/sub0/c13 ),
    .f(\trig_node/trigger_node_int_0/n141 [14:13]),
    .fco(\trig_node/trigger_node_int_0/sub0/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/sub0/u0|trig_node/trigger_node_int_0/sub0/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/sub0/u15_al_u3569  (
    .a({open_n44830,control_21}),
    .b({open_n44831,1'b0}),
    .fci(\trig_node/trigger_node_int_0/sub0/c15 ),
    .f({open_n44850,\trig_node/trigger_node_int_0/n141 [15]}));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/sub0/u0|trig_node/trigger_node_int_0/sub0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/sub0/u2|trig_node/trigger_node_int_0/sub0/u1  (
    .a({control_8,control_7}),
    .b(2'b01),
    .fci(\trig_node/trigger_node_int_0/sub0/c1 ),
    .f(\trig_node/trigger_node_int_0/n141 [2:1]),
    .fco(\trig_node/trigger_node_int_0/sub0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/sub0/u0|trig_node/trigger_node_int_0/sub0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/sub0/u4|trig_node/trigger_node_int_0/sub0/u3  (
    .a({control_10,control_9}),
    .b(2'b01),
    .fci(\trig_node/trigger_node_int_0/sub0/c3 ),
    .f(\trig_node/trigger_node_int_0/n141 [4:3]),
    .fco(\trig_node/trigger_node_int_0/sub0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/sub0/u0|trig_node/trigger_node_int_0/sub0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/sub0/u6|trig_node/trigger_node_int_0/sub0/u5  (
    .a({control_12,control_11}),
    .b(2'b01),
    .fci(\trig_node/trigger_node_int_0/sub0/c5 ),
    .f(\trig_node/trigger_node_int_0/n141 [6:5]),
    .fco(\trig_node/trigger_node_int_0/sub0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("trig_node/trigger_node_int_0/sub0/u0|trig_node/trigger_node_int_0/sub0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \trig_node/trigger_node_int_0/sub0/u8|trig_node/trigger_node_int_0/sub0/u7  (
    .a({control_14,control_13}),
    .b(2'b00),
    .fci(\trig_node/trigger_node_int_0/sub0/c7 ),
    .f(\trig_node/trigger_node_int_0/n141 [8:7]),
    .fco(\trig_node/trigger_node_int_0/sub0/c9 ));
  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/trig_rstn_sync0_reg|trig_node/trigger_node_int_0/trig_rstn_sync_reg  (
    .clk(clock_pad),
    .mi({control_0,\trig_node/trigger_node_int_0/trig_rstn_sync0 }),
    .q({\trig_node/trigger_node_int_0/trig_rstn_sync0 ,\trig_node/trigger_node_int_0/trig_rstn_sync }));  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/trig_rstn_sync0_reg|trig_node/trigger_node_int_0/trig_rstn_sync_reg_placeOpt_1  (
    .clk(clock_pad),
    .mi({control_0,\trig_node/trigger_node_int_0/trig_rstn_sync0 }),
    .q({open_n45002,\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_1 }));  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/trig_rstn_sync0_reg|trig_node/trigger_node_int_0/trig_rstn_sync_reg_placeOpt_10  (
    .clk(clock_pad),
    .mi({control_0,\trig_node/trigger_node_int_0/trig_rstn_sync0 }),
    .q({open_n45032,\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_10 }));  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/trig_rstn_sync0_reg|trig_node/trigger_node_int_0/trig_rstn_sync_reg_placeOpt_2  (
    .clk(clock_pad),
    .mi({control_0,\trig_node/trigger_node_int_0/trig_rstn_sync0 }),
    .q({open_n45062,\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_2 }));  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/trig_rstn_sync0_reg|trig_node/trigger_node_int_0/trig_rstn_sync_reg_placeOpt_3  (
    .clk(clock_pad),
    .mi({control_0,\trig_node/trigger_node_int_0/trig_rstn_sync0 }),
    .q({open_n45092,\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_3 }));  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/trig_rstn_sync0_reg|trig_node/trigger_node_int_0/trig_rstn_sync_reg_placeOpt_4  (
    .clk(clock_pad),
    .mi({control_0,\trig_node/trigger_node_int_0/trig_rstn_sync0 }),
    .q({open_n45122,\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_4 }));  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/trig_rstn_sync0_reg|trig_node/trigger_node_int_0/trig_rstn_sync_reg_placeOpt_5  (
    .clk(clock_pad),
    .mi({control_0,\trig_node/trigger_node_int_0/trig_rstn_sync0 }),
    .q({open_n45152,\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_5 }));  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/trig_rstn_sync0_reg|trig_node/trigger_node_int_0/trig_rstn_sync_reg_placeOpt_6  (
    .clk(clock_pad),
    .mi({control_0,\trig_node/trigger_node_int_0/trig_rstn_sync0 }),
    .q({open_n45182,\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_6 }));  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/trig_rstn_sync0_reg|trig_node/trigger_node_int_0/trig_rstn_sync_reg_placeOpt_7  (
    .clk(clock_pad),
    .mi({control_0,\trig_node/trigger_node_int_0/trig_rstn_sync0 }),
    .q({open_n45212,\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_7 }));  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/trig_rstn_sync0_reg|trig_node/trigger_node_int_0/trig_rstn_sync_reg_placeOpt_8  (
    .clk(clock_pad),
    .mi({control_0,\trig_node/trigger_node_int_0/trig_rstn_sync0 }),
    .q({open_n45242,\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_8 }));  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_LSLICE #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \trig_node/trigger_node_int_0/trig_rstn_sync0_reg|trig_node/trigger_node_int_0/trig_rstn_sync_reg_placeOpt_9  (
    .clk(clock_pad),
    .mi({control_0,\trig_node/trigger_node_int_0/trig_rstn_sync0 }),
    .q({open_n45272,\trig_node/trigger_node_int_0/trig_rstn_sync_placeOpt_9 }));  // D:/td/td/cw\trigger_node.v(47)
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1/u0|u1/ucin  (
    .a({\t/memstraddress [2],1'b0}),
    .b({1'b1,open_n45273}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .mi({open_n45288,\t/memstraddress [2]}),
    .sr(rst_pad),
    .f({n4[0],open_n45289}),
    .fco(\u1/c1 ),
    .q({open_n45292,\t/a/ID_memstraddr [2]}));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u10|u1/u9  (
    .a(\t/memstraddress [12:11]),
    .b(2'b00),
    .fci(\u1/c9 ),
    .f(n4[10:9]),
    .fco(\u1/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u12|u1/u11  (
    .a(\t/memstraddress [14:13]),
    .b(2'b00),
    .fci(\u1/c11 ),
    .f(n4[12:11]),
    .fco(\u1/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u14|u1/u13  (
    .a(\t/memstraddress [16:15]),
    .b(2'b00),
    .fci(\u1/c13 ),
    .f(n4[14:13]),
    .fco(\u1/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u16|u1/u15  (
    .a(\t/memstraddress [18:17]),
    .b(2'b00),
    .fci(\u1/c15 ),
    .f(n4[16:15]),
    .fco(\u1/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u18|u1/u17  (
    .a(\t/memstraddress [20:19]),
    .b(2'b00),
    .fci(\u1/c17 ),
    .f(n4[18:17]),
    .fco(\u1/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u20|u1/u19  (
    .a(\t/memstraddress [22:21]),
    .b(2'b00),
    .fci(\u1/c19 ),
    .f(n4[20:19]),
    .fco(\u1/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u22|u1/u21  (
    .a(\t/memstraddress [24:23]),
    .b(2'b00),
    .fci(\u1/c21 ),
    .f(n4[22:21]),
    .fco(\u1/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u24|u1/u23  (
    .a(\t/memstraddress [26:25]),
    .b(2'b00),
    .fci(\u1/c23 ),
    .f(n4[24:23]),
    .fco(\u1/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u26|u1/u25  (
    .a(\t/memstraddress [28:27]),
    .b(2'b00),
    .fci(\u1/c25 ),
    .f(n4[26:25]),
    .fco(\u1/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u28|u1/u27  (
    .a(\t/memstraddress [30:29]),
    .b(2'b00),
    .fci(\u1/c27 ),
    .f(n4[28:27]),
    .fco(\u1/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u29_al_u2978  (
    .a({open_n45513,\t/memstraddress [31]}),
    .b({open_n45514,1'b0}),
    .fci(\u1/c29 ),
    .f({open_n45533,n4[29]}));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u2|u1/u1  (
    .a(\t/memstraddress [4:3]),
    .b(2'b00),
    .fci(\u1/c1 ),
    .f(n4[2:1]),
    .fco(\u1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u4|u1/u3  (
    .a(\t/memstraddress [6:5]),
    .b(2'b00),
    .fci(\u1/c3 ),
    .f(n4[4:3]),
    .fco(\u1/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u6|u1/u5  (
    .a(\t/memstraddress [8:7]),
    .b(2'b00),
    .fci(\u1/c5 ),
    .f(n4[6:5]),
    .fco(\u1/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u8|u1/u7  (
    .a(\t/memstraddress [10:9]),
    .b(2'b00),
    .fci(\u1/c7 ),
    .f(n4[8:7]),
    .fco(\u1/c9 ));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u11_al_u2964  (
    .a({\t/a/ID_jump_addr [14],\t/a/ID_jump_addr [12]}),
    .b({\t/a/ID_jump_addr [15],\t/a/ID_jump_addr [13]}),
    .c(2'b00),
    .d({n4[12],n4[10]}),
    .e({n4[13],n4[11]}),
    .fci(\u3/c11 ),
    .f({n8[13],n8[11]}),
    .fco(\u3/c15 ),
    .fx({n8[14],n8[12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u15_al_u2965  (
    .a({\t/a/ID_jump_addr [18],\t/a/ID_jump_addr [16]}),
    .b({\t/a/ID_jump_addr [19],\t/a/ID_jump_addr [17]}),
    .c(2'b00),
    .d({n4[16],n4[14]}),
    .e({n4[17],n4[15]}),
    .fci(\u3/c15 ),
    .f({n8[17],n8[15]}),
    .fco(\u3/c19 ),
    .fx({n8[18],n8[16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u19_al_u2966  (
    .a({\t/a/ID_jump_addr [22],\t/a/ID_jump_addr [20]}),
    .b({\t/a/ID_jump_addr [23],\t/a/ID_jump_addr [21]}),
    .c(2'b00),
    .d({n4[20],n4[18]}),
    .e({n4[21],n4[19]}),
    .fci(\u3/c19 ),
    .f({n8[21],n8[19]}),
    .fco(\u3/c23 ),
    .fx({n8[22],n8[20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u23_al_u2967  (
    .a({\t/a/ID_jump_addr [26],\t/a/ID_jump_addr [24]}),
    .b({\t/a/ID_jump_addr [27],\t/a/ID_jump_addr [25]}),
    .c(2'b00),
    .d({n4[24],n4[22]}),
    .e({n4[25],n4[23]}),
    .fci(\u3/c23 ),
    .f({n8[25],n8[23]}),
    .fco(\u3/c27 ),
    .fx({n8[26],n8[24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u27_al_u2968  (
    .a({\t/a/ID_jump_addr [30],\t/a/ID_jump_addr [28]}),
    .b({\t/a/ID_jump_addr [31],\t/a/ID_jump_addr [29]}),
    .c(2'b00),
    .d({n4[28],n4[26]}),
    .e({n4[29],n4[27]}),
    .fci(\u3/c27 ),
    .f({n8[29],n8[27]}),
    .fx({n8[30],n8[28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u3_al_u2962  (
    .a({\t/a/ID_jump_addr [6],\t/a/ID_jump_addr [4]}),
    .b({\t/a/ID_jump_addr [7],\t/a/ID_jump_addr [5]}),
    .c(2'b00),
    .d({n4[4],n4[2]}),
    .e({n4[5],n4[3]}),
    .fci(\u3/c3 ),
    .f({n8[5],n8[3]}),
    .fco(\u3/c7 ),
    .fx({n8[6],n8[4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u7_al_u2963  (
    .a({\t/a/ID_jump_addr [10],\t/a/ID_jump_addr [8]}),
    .b({\t/a/ID_jump_addr [11],\t/a/ID_jump_addr [9]}),
    .c(2'b00),
    .d({n4[8],n4[6]}),
    .e({n4[9],n4[7]}),
    .fci(\u3/c7 ),
    .f({n8[9],n8[7]}),
    .fco(\u3/c11 ),
    .fx({n8[10],n8[8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u3/ucin_al_u2961  (
    .a({\t/a/ID_jump_addr [2],1'b0}),
    .b({\t/a/ID_jump_addr [3],\t/a/ID_jump_addr [1]}),
    .c(2'b00),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({n4[0],1'b1}),
    .e({n4[1],\t/memstraddress [1]}),
    .mi({open_n45755,\t/memstraddress [1]}),
    .sr(rst_pad),
    .f({n8[1],open_n45767}),
    .fco(\u3/c3 ),
    .fx({n8[2],n8[0]}),
    .q({open_n45768,\t/a/ID_memstraddr [1]}));

endmodule 

