// Verilog netlist created by TD v4.3.815
// Fri Mar 22 13:53:44 2019

`timescale 1ns / 1ps
module __top  // __top.v(3)
  (
  clock,
  rst,
  led
  );

  input clock;  // __top.v(4)
  input rst;  // __top.v(3)
  output led;  // __top.v(5)

  wire [31:0] addr;  // __top.v(17)
  wire [31:0] i_data;  // __top.v(15)
  wire [3:0] \m/dram_c0_di ;
  wire [3:0] \m/dram_c0_waddr ;
  wire [3:0] \m/dram_c1_di ;
  wire [3:0] \m/dram_c1_waddr ;
  wire [3:0] \m/dram_c2_di ;
  wire [3:0] \m/dram_c2_waddr ;
  wire [3:0] \m/dram_c3_di ;
  wire [3:0] \m/dram_c3_waddr ;
  wire [3:0] \m/dram_c4_di ;
  wire [3:0] \m/dram_c4_waddr ;
  wire [3:0] \m/dram_c5_di ;
  wire [3:0] \m/dram_c5_waddr ;
  wire [3:0] \m/dram_c6_di ;
  wire [3:0] \m/dram_c6_waddr ;
  wire [3:0] \m/dram_c7_di ;
  wire [3:0] \m/dram_c7_waddr ;
  wire [3:0] n2;
  wire [3:0] n3;
  wire [29:0] n4;
  wire [30:0] n8;
  wire [31:0] o_data;  // __top.v(16)
  wire [31:0] \t/a/EX_A ;  // cpu.v(47)
  wire [31:0] \t/a/EX_B ;  // cpu.v(48)
  wire [2:0] \t/a/EX_fun3 ;  // cpu.v(49)
  wire [6:0] \t/a/EX_fun7 ;  // cpu.v(41)
  wire [31:0] \t/a/EX_memstraddr ;  // cpu.v(38)
  wire [6:0] \t/a/EX_op ;  // cpu.v(42)
  wire [3:0] \t/a/EX_operation ;  // cpu.v(46)
  wire [4:0] \t/a/EX_rd ;  // cpu.v(45)
  wire [31:0] \t/a/EX_regdat1 ;  // cpu.v(39)
  wire [31:0] \t/a/EX_regdat2 ;  // cpu.v(40)
  wire [4:0] \t/a/EX_rs1 ;  // cpu.v(43)
  wire [4:0] \t/a/EX_rs2 ;  // cpu.v(44)
  wire [2:0] \t/a/ID_fun3 ;  // cpu.v(21)
  wire [6:0] \t/a/ID_fun7 ;  // cpu.v(22)
  wire [31:0] \t/a/ID_jump_addr ;  // cpu.v(28)
  wire [31:0] \t/a/ID_jump_regdat1 ;  // cpu.v(29)
  wire [31:0] \t/a/ID_jump_regdat2 ;  // cpu.v(30)
  wire [31:0] \t/a/ID_memstraddr ;  // cpu.v(26)
  wire [6:0] \t/a/ID_op ;  // cpu.v(20)
  wire [4:0] \t/a/ID_rd ;  // cpu.v(23)
  wire [31:0] \t/a/ID_read_dat1 ;  // cpu.v(36)
  wire [31:0] \t/a/ID_read_dat2 ;  // cpu.v(37)
  wire [4:0] \t/a/ID_rs1 ;  // cpu.v(24)
  wire [4:0] \t/a/ID_rs2 ;  // cpu.v(25)
  wire [31:0] \t/a/IF_skip_addr ;  // cpu.v(17)
  wire [31:0] \t/a/MEM_aludat ;  // cpu.v(54)
  wire [2:0] \t/a/MEM_fun3 ;  // cpu.v(58)
  wire [6:0] \t/a/MEM_op ;  // cpu.v(55)
  wire [4:0] \t/a/MEM_rd ;  // cpu.v(56)
  wire [31:0] \t/a/MEM_regdat2 ;  // cpu.v(57)
  wire [6:0] \t/a/WB_op ;  // cpu.v(71)
  wire [4:0] \t/a/WB_rd ;  // cpu.v(70)
  wire  \t/a/alu/mux0_b1/B1_0 ;
  wire  \t/a/alu/mux0_b2/B1_0 ;
  wire  \t/a/alu/mux0_b3/B1_0 ;
  wire  \t/a/alu/mux0_b5/B1_0 ;
  wire  \t/a/alu/mux0_b6/B1_0 ;
  wire [31:0] \t/a/alu/n5 ;
  wire [31:0] \t/a/alu/n6 ;
  wire [1:0] \t/a/alu_A_select ;  // cpu.v(33)
  wire [1:0] \t/a/alu_B_select ;  // cpu.v(34)
  wire [31:0] \t/a/aludat ;  // cpu.v(52)
  wire  \t/a/aluin/sel0_b0/B0 ;
  wire  \t/a/aluin/sel0_b1/B0 ;
  wire  \t/a/aluin/sel0_b10/B0 ;
  wire  \t/a/aluin/sel0_b11/B0 ;
  wire  \t/a/aluin/sel0_b12/B0 ;
  wire  \t/a/aluin/sel0_b13/B0 ;
  wire  \t/a/aluin/sel0_b14/B0 ;
  wire  \t/a/aluin/sel0_b15/B0 ;
  wire  \t/a/aluin/sel0_b16/B0 ;
  wire  \t/a/aluin/sel0_b17/B0 ;
  wire  \t/a/aluin/sel0_b18/B0 ;
  wire  \t/a/aluin/sel0_b19/B0 ;
  wire  \t/a/aluin/sel0_b2/B0 ;
  wire  \t/a/aluin/sel0_b20/B0 ;
  wire  \t/a/aluin/sel0_b21/B0 ;
  wire  \t/a/aluin/sel0_b22/B0 ;
  wire  \t/a/aluin/sel0_b23/B0 ;
  wire  \t/a/aluin/sel0_b24/B0 ;
  wire  \t/a/aluin/sel0_b25/B0 ;
  wire  \t/a/aluin/sel0_b26/B0 ;
  wire  \t/a/aluin/sel0_b27/B0 ;
  wire  \t/a/aluin/sel0_b28/B0 ;
  wire  \t/a/aluin/sel0_b29/B0 ;
  wire  \t/a/aluin/sel0_b3/B0 ;
  wire  \t/a/aluin/sel0_b30/B0 ;
  wire  \t/a/aluin/sel0_b31/B0 ;
  wire  \t/a/aluin/sel0_b4/B0 ;
  wire  \t/a/aluin/sel0_b5/B0 ;
  wire  \t/a/aluin/sel0_b6/B0 ;
  wire  \t/a/aluin/sel0_b7/B0 ;
  wire  \t/a/aluin/sel0_b8/B0 ;
  wire  \t/a/aluin/sel0_b9/B0 ;
  wire  \t/a/aluin/sel1_b10/B9 ;
  wire  \t/a/aluin/sel1_b11/B9 ;
  wire  \t/a/aluin/sel1_b12/B9 ;
  wire  \t/a/aluin/sel1_b13/B9 ;
  wire  \t/a/aluin/sel1_b14/B9 ;
  wire  \t/a/aluin/sel1_b15/B9 ;
  wire  \t/a/aluin/sel1_b16/B9 ;
  wire  \t/a/aluin/sel1_b17/B9 ;
  wire  \t/a/aluin/sel1_b18/B9 ;
  wire  \t/a/aluin/sel1_b19/B9 ;
  wire  \t/a/aluin/sel1_b20/B9 ;
  wire  \t/a/aluin/sel1_b21/B9 ;
  wire  \t/a/aluin/sel1_b22/B9 ;
  wire  \t/a/aluin/sel1_b23/B9 ;
  wire  \t/a/aluin/sel1_b24/B9 ;
  wire  \t/a/aluin/sel1_b25/B9 ;
  wire  \t/a/aluin/sel1_b26/B9 ;
  wire  \t/a/aluin/sel1_b27/B9 ;
  wire  \t/a/aluin/sel1_b28/B9 ;
  wire  \t/a/aluin/sel1_b29/B9 ;
  wire  \t/a/aluin/sel1_b30/B9 ;
  wire  \t/a/aluin/sel1_b31/B9 ;
  wire  \t/a/aluin/sel1_b5/B9 ;
  wire  \t/a/aluin/sel1_b6/B9 ;
  wire  \t/a/aluin/sel1_b7/B9 ;
  wire  \t/a/aluin/sel1_b8/B9 ;
  wire  \t/a/aluin/sel1_b9/B9 ;
  wire [31:0] \t/a/condition/n3 ;
  wire [31:0] \t/a/condition/n5 ;
  wire  \t/a/condition/sel0_b12/B1 ;
  wire  \t/a/condition/sel1/B2 ;
  wire [31:0] \t/a/instr/n12 ;
  wire [29:0] \t/a/instr/n16 ;
  wire  \t/a/mux4_b7/B0_0 ;
  wire [31:0] \t/a/reg_writedat ;  // cpu.v(68)
  wire [31:0] \t/a/regfile/n46 ;
  wire [31:0] \t/a/regfile/regfile$0$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$1$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$10$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$11$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$12$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$13$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$14$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$15$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$16$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$17$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$18$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$19$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$2$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$20$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$21$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$22$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$23$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$24$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$25$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$26$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$27$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$28$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$29$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$3$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$30$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$31$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$4$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$5$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$6$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$7$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$8$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$9$ ;  // register.v(5)
  wire [31:0] \t/busarbitration/instruction ;  // io.v(35)
  wire [31:0] \t/memstraddress ;  // top2.v(17)
  wire _al_u1000_o;
  wire _al_u1001_o;
  wire _al_u1002_o;
  wire _al_u1003_o;
  wire _al_u1004_o;
  wire _al_u1043_o;
  wire _al_u1044_o;
  wire _al_u1045_o;
  wire _al_u1046_o;
  wire _al_u1047_o;
  wire _al_u1049_o;
  wire _al_u1050_o;
  wire _al_u1051_o;
  wire _al_u1052_o;
  wire _al_u1053_o;
  wire _al_u1054_o;
  wire _al_u1055_o;
  wire _al_u1056_o;
  wire _al_u1057_o;
  wire _al_u1058_o;
  wire _al_u1059_o;
  wire _al_u1060_o;
  wire _al_u1061_o;
  wire _al_u1062_o;
  wire _al_u1063_o;
  wire _al_u1064_o;
  wire _al_u1065_o;
  wire _al_u1066_o;
  wire _al_u1067_o;
  wire _al_u1068_o;
  wire _al_u1069_o;
  wire _al_u1071_o;
  wire _al_u1072_o;
  wire _al_u1073_o;
  wire _al_u1074_o;
  wire _al_u1075_o;
  wire _al_u1076_o;
  wire _al_u1077_o;
  wire _al_u1078_o;
  wire _al_u1079_o;
  wire _al_u1080_o;
  wire _al_u1081_o;
  wire _al_u1082_o;
  wire _al_u1083_o;
  wire _al_u1084_o;
  wire _al_u1085_o;
  wire _al_u1086_o;
  wire _al_u1087_o;
  wire _al_u1088_o;
  wire _al_u1089_o;
  wire _al_u1090_o;
  wire _al_u1092_o;
  wire _al_u1093_o;
  wire _al_u1094_o;
  wire _al_u1095_o;
  wire _al_u1096_o;
  wire _al_u1097_o;
  wire _al_u1098_o;
  wire _al_u1099_o;
  wire _al_u1100_o;
  wire _al_u1101_o;
  wire _al_u1102_o;
  wire _al_u1103_o;
  wire _al_u1104_o;
  wire _al_u1105_o;
  wire _al_u1106_o;
  wire _al_u1107_o;
  wire _al_u1108_o;
  wire _al_u1109_o;
  wire _al_u1110_o;
  wire _al_u1111_o;
  wire _al_u1113_o;
  wire _al_u1114_o;
  wire _al_u1115_o;
  wire _al_u1116_o;
  wire _al_u1117_o;
  wire _al_u1118_o;
  wire _al_u1119_o;
  wire _al_u1120_o;
  wire _al_u1121_o;
  wire _al_u1122_o;
  wire _al_u1123_o;
  wire _al_u1124_o;
  wire _al_u1125_o;
  wire _al_u1126_o;
  wire _al_u1127_o;
  wire _al_u1128_o;
  wire _al_u1129_o;
  wire _al_u1130_o;
  wire _al_u1131_o;
  wire _al_u1132_o;
  wire _al_u1134_o;
  wire _al_u1135_o;
  wire _al_u1136_o;
  wire _al_u1137_o;
  wire _al_u1138_o;
  wire _al_u1139_o;
  wire _al_u1140_o;
  wire _al_u1141_o;
  wire _al_u1142_o;
  wire _al_u1143_o;
  wire _al_u1144_o;
  wire _al_u1145_o;
  wire _al_u1146_o;
  wire _al_u1147_o;
  wire _al_u1148_o;
  wire _al_u1149_o;
  wire _al_u1150_o;
  wire _al_u1151_o;
  wire _al_u1152_o;
  wire _al_u1153_o;
  wire _al_u1155_o;
  wire _al_u1156_o;
  wire _al_u1157_o;
  wire _al_u1158_o;
  wire _al_u1159_o;
  wire _al_u1160_o;
  wire _al_u1161_o;
  wire _al_u1162_o;
  wire _al_u1163_o;
  wire _al_u1164_o;
  wire _al_u1165_o;
  wire _al_u1166_o;
  wire _al_u1167_o;
  wire _al_u1168_o;
  wire _al_u1169_o;
  wire _al_u1170_o;
  wire _al_u1171_o;
  wire _al_u1172_o;
  wire _al_u1173_o;
  wire _al_u1174_o;
  wire _al_u1176_o;
  wire _al_u1177_o;
  wire _al_u1178_o;
  wire _al_u1179_o;
  wire _al_u1180_o;
  wire _al_u1181_o;
  wire _al_u1182_o;
  wire _al_u1183_o;
  wire _al_u1184_o;
  wire _al_u1185_o;
  wire _al_u1186_o;
  wire _al_u1187_o;
  wire _al_u1188_o;
  wire _al_u1189_o;
  wire _al_u1190_o;
  wire _al_u1191_o;
  wire _al_u1192_o;
  wire _al_u1193_o;
  wire _al_u1194_o;
  wire _al_u1195_o;
  wire _al_u1197_o;
  wire _al_u1198_o;
  wire _al_u1199_o;
  wire _al_u1200_o;
  wire _al_u1201_o;
  wire _al_u1202_o;
  wire _al_u1203_o;
  wire _al_u1204_o;
  wire _al_u1205_o;
  wire _al_u1206_o;
  wire _al_u1207_o;
  wire _al_u1208_o;
  wire _al_u1209_o;
  wire _al_u1210_o;
  wire _al_u1211_o;
  wire _al_u1212_o;
  wire _al_u1213_o;
  wire _al_u1214_o;
  wire _al_u1215_o;
  wire _al_u1216_o;
  wire _al_u1218_o;
  wire _al_u1219_o;
  wire _al_u1220_o;
  wire _al_u1221_o;
  wire _al_u1222_o;
  wire _al_u1223_o;
  wire _al_u1224_o;
  wire _al_u1225_o;
  wire _al_u1226_o;
  wire _al_u1227_o;
  wire _al_u1228_o;
  wire _al_u1229_o;
  wire _al_u1230_o;
  wire _al_u1231_o;
  wire _al_u1232_o;
  wire _al_u1233_o;
  wire _al_u1234_o;
  wire _al_u1235_o;
  wire _al_u1236_o;
  wire _al_u1237_o;
  wire _al_u1239_o;
  wire _al_u1240_o;
  wire _al_u1241_o;
  wire _al_u1242_o;
  wire _al_u1243_o;
  wire _al_u1244_o;
  wire _al_u1245_o;
  wire _al_u1246_o;
  wire _al_u1247_o;
  wire _al_u1248_o;
  wire _al_u1249_o;
  wire _al_u1250_o;
  wire _al_u1251_o;
  wire _al_u1252_o;
  wire _al_u1253_o;
  wire _al_u1254_o;
  wire _al_u1255_o;
  wire _al_u1256_o;
  wire _al_u1257_o;
  wire _al_u1258_o;
  wire _al_u1260_o;
  wire _al_u1261_o;
  wire _al_u1262_o;
  wire _al_u1263_o;
  wire _al_u1264_o;
  wire _al_u1265_o;
  wire _al_u1266_o;
  wire _al_u1267_o;
  wire _al_u1268_o;
  wire _al_u1269_o;
  wire _al_u1270_o;
  wire _al_u1271_o;
  wire _al_u1272_o;
  wire _al_u1273_o;
  wire _al_u1274_o;
  wire _al_u1275_o;
  wire _al_u1276_o;
  wire _al_u1277_o;
  wire _al_u1278_o;
  wire _al_u1279_o;
  wire _al_u1281_o;
  wire _al_u1282_o;
  wire _al_u1283_o;
  wire _al_u1284_o;
  wire _al_u1285_o;
  wire _al_u1286_o;
  wire _al_u1287_o;
  wire _al_u1288_o;
  wire _al_u1289_o;
  wire _al_u1290_o;
  wire _al_u1291_o;
  wire _al_u1292_o;
  wire _al_u1293_o;
  wire _al_u1294_o;
  wire _al_u1295_o;
  wire _al_u1296_o;
  wire _al_u1297_o;
  wire _al_u1298_o;
  wire _al_u1299_o;
  wire _al_u1300_o;
  wire _al_u1302_o;
  wire _al_u1303_o;
  wire _al_u1304_o;
  wire _al_u1305_o;
  wire _al_u1306_o;
  wire _al_u1307_o;
  wire _al_u1308_o;
  wire _al_u1309_o;
  wire _al_u1310_o;
  wire _al_u1311_o;
  wire _al_u1312_o;
  wire _al_u1313_o;
  wire _al_u1314_o;
  wire _al_u1315_o;
  wire _al_u1316_o;
  wire _al_u1317_o;
  wire _al_u1318_o;
  wire _al_u1319_o;
  wire _al_u1320_o;
  wire _al_u1321_o;
  wire _al_u1323_o;
  wire _al_u1324_o;
  wire _al_u1325_o;
  wire _al_u1326_o;
  wire _al_u1327_o;
  wire _al_u1328_o;
  wire _al_u1329_o;
  wire _al_u1330_o;
  wire _al_u1331_o;
  wire _al_u1332_o;
  wire _al_u1333_o;
  wire _al_u1334_o;
  wire _al_u1335_o;
  wire _al_u1336_o;
  wire _al_u1337_o;
  wire _al_u1338_o;
  wire _al_u1339_o;
  wire _al_u1340_o;
  wire _al_u1341_o;
  wire _al_u1342_o;
  wire _al_u1344_o;
  wire _al_u1345_o;
  wire _al_u1346_o;
  wire _al_u1347_o;
  wire _al_u1348_o;
  wire _al_u1349_o;
  wire _al_u1350_o;
  wire _al_u1351_o;
  wire _al_u1352_o;
  wire _al_u1353_o;
  wire _al_u1354_o;
  wire _al_u1355_o;
  wire _al_u1356_o;
  wire _al_u1357_o;
  wire _al_u1358_o;
  wire _al_u1359_o;
  wire _al_u1360_o;
  wire _al_u1361_o;
  wire _al_u1362_o;
  wire _al_u1363_o;
  wire _al_u1365_o;
  wire _al_u1366_o;
  wire _al_u1367_o;
  wire _al_u1368_o;
  wire _al_u1369_o;
  wire _al_u1370_o;
  wire _al_u1371_o;
  wire _al_u1372_o;
  wire _al_u1373_o;
  wire _al_u1374_o;
  wire _al_u1375_o;
  wire _al_u1376_o;
  wire _al_u1377_o;
  wire _al_u1378_o;
  wire _al_u1379_o;
  wire _al_u1380_o;
  wire _al_u1381_o;
  wire _al_u1382_o;
  wire _al_u1383_o;
  wire _al_u1384_o;
  wire _al_u1386_o;
  wire _al_u1387_o;
  wire _al_u1388_o;
  wire _al_u1389_o;
  wire _al_u1390_o;
  wire _al_u1391_o;
  wire _al_u1392_o;
  wire _al_u1393_o;
  wire _al_u1394_o;
  wire _al_u1395_o;
  wire _al_u1396_o;
  wire _al_u1397_o;
  wire _al_u1398_o;
  wire _al_u1399_o;
  wire _al_u1400_o;
  wire _al_u1401_o;
  wire _al_u1402_o;
  wire _al_u1403_o;
  wire _al_u1404_o;
  wire _al_u1405_o;
  wire _al_u1407_o;
  wire _al_u1408_o;
  wire _al_u1409_o;
  wire _al_u1410_o;
  wire _al_u1411_o;
  wire _al_u1412_o;
  wire _al_u1413_o;
  wire _al_u1414_o;
  wire _al_u1415_o;
  wire _al_u1416_o;
  wire _al_u1417_o;
  wire _al_u1418_o;
  wire _al_u1419_o;
  wire _al_u1420_o;
  wire _al_u1421_o;
  wire _al_u1422_o;
  wire _al_u1423_o;
  wire _al_u1424_o;
  wire _al_u1425_o;
  wire _al_u1426_o;
  wire _al_u1428_o;
  wire _al_u1429_o;
  wire _al_u1430_o;
  wire _al_u1431_o;
  wire _al_u1432_o;
  wire _al_u1433_o;
  wire _al_u1434_o;
  wire _al_u1435_o;
  wire _al_u1436_o;
  wire _al_u1437_o;
  wire _al_u1438_o;
  wire _al_u1439_o;
  wire _al_u1440_o;
  wire _al_u1441_o;
  wire _al_u1442_o;
  wire _al_u1443_o;
  wire _al_u1444_o;
  wire _al_u1445_o;
  wire _al_u1446_o;
  wire _al_u1447_o;
  wire _al_u1449_o;
  wire _al_u1450_o;
  wire _al_u1451_o;
  wire _al_u1452_o;
  wire _al_u1453_o;
  wire _al_u1454_o;
  wire _al_u1455_o;
  wire _al_u1456_o;
  wire _al_u1457_o;
  wire _al_u1458_o;
  wire _al_u1459_o;
  wire _al_u1460_o;
  wire _al_u1461_o;
  wire _al_u1462_o;
  wire _al_u1463_o;
  wire _al_u1464_o;
  wire _al_u1465_o;
  wire _al_u1466_o;
  wire _al_u1467_o;
  wire _al_u1468_o;
  wire _al_u1470_o;
  wire _al_u1471_o;
  wire _al_u1472_o;
  wire _al_u1473_o;
  wire _al_u1474_o;
  wire _al_u1475_o;
  wire _al_u1476_o;
  wire _al_u1477_o;
  wire _al_u1478_o;
  wire _al_u1479_o;
  wire _al_u1480_o;
  wire _al_u1481_o;
  wire _al_u1482_o;
  wire _al_u1483_o;
  wire _al_u1484_o;
  wire _al_u1485_o;
  wire _al_u1486_o;
  wire _al_u1487_o;
  wire _al_u1488_o;
  wire _al_u1489_o;
  wire _al_u1491_o;
  wire _al_u1492_o;
  wire _al_u1493_o;
  wire _al_u1494_o;
  wire _al_u1495_o;
  wire _al_u1496_o;
  wire _al_u1497_o;
  wire _al_u1498_o;
  wire _al_u1499_o;
  wire _al_u1500_o;
  wire _al_u1501_o;
  wire _al_u1502_o;
  wire _al_u1503_o;
  wire _al_u1504_o;
  wire _al_u1505_o;
  wire _al_u1506_o;
  wire _al_u1507_o;
  wire _al_u1508_o;
  wire _al_u1509_o;
  wire _al_u1510_o;
  wire _al_u1512_o;
  wire _al_u1513_o;
  wire _al_u1514_o;
  wire _al_u1515_o;
  wire _al_u1516_o;
  wire _al_u1517_o;
  wire _al_u1518_o;
  wire _al_u1519_o;
  wire _al_u1520_o;
  wire _al_u1521_o;
  wire _al_u1522_o;
  wire _al_u1523_o;
  wire _al_u1524_o;
  wire _al_u1525_o;
  wire _al_u1526_o;
  wire _al_u1527_o;
  wire _al_u1528_o;
  wire _al_u1529_o;
  wire _al_u1530_o;
  wire _al_u1531_o;
  wire _al_u1533_o;
  wire _al_u1534_o;
  wire _al_u1535_o;
  wire _al_u1536_o;
  wire _al_u1537_o;
  wire _al_u1538_o;
  wire _al_u1539_o;
  wire _al_u1540_o;
  wire _al_u1541_o;
  wire _al_u1542_o;
  wire _al_u1543_o;
  wire _al_u1544_o;
  wire _al_u1545_o;
  wire _al_u1546_o;
  wire _al_u1547_o;
  wire _al_u1548_o;
  wire _al_u1549_o;
  wire _al_u1550_o;
  wire _al_u1551_o;
  wire _al_u1552_o;
  wire _al_u1554_o;
  wire _al_u1555_o;
  wire _al_u1556_o;
  wire _al_u1557_o;
  wire _al_u1558_o;
  wire _al_u1559_o;
  wire _al_u1560_o;
  wire _al_u1561_o;
  wire _al_u1562_o;
  wire _al_u1563_o;
  wire _al_u1564_o;
  wire _al_u1565_o;
  wire _al_u1566_o;
  wire _al_u1567_o;
  wire _al_u1568_o;
  wire _al_u1569_o;
  wire _al_u1570_o;
  wire _al_u1571_o;
  wire _al_u1572_o;
  wire _al_u1573_o;
  wire _al_u1575_o;
  wire _al_u1576_o;
  wire _al_u1577_o;
  wire _al_u1578_o;
  wire _al_u1579_o;
  wire _al_u1580_o;
  wire _al_u1581_o;
  wire _al_u1582_o;
  wire _al_u1583_o;
  wire _al_u1584_o;
  wire _al_u1585_o;
  wire _al_u1586_o;
  wire _al_u1587_o;
  wire _al_u1588_o;
  wire _al_u1589_o;
  wire _al_u1590_o;
  wire _al_u1591_o;
  wire _al_u1592_o;
  wire _al_u1593_o;
  wire _al_u1594_o;
  wire _al_u1596_o;
  wire _al_u1597_o;
  wire _al_u1598_o;
  wire _al_u1599_o;
  wire _al_u1600_o;
  wire _al_u1601_o;
  wire _al_u1602_o;
  wire _al_u1603_o;
  wire _al_u1604_o;
  wire _al_u1605_o;
  wire _al_u1606_o;
  wire _al_u1607_o;
  wire _al_u1608_o;
  wire _al_u1609_o;
  wire _al_u1610_o;
  wire _al_u1611_o;
  wire _al_u1612_o;
  wire _al_u1613_o;
  wire _al_u1614_o;
  wire _al_u1615_o;
  wire _al_u1617_o;
  wire _al_u1618_o;
  wire _al_u1619_o;
  wire _al_u1620_o;
  wire _al_u1621_o;
  wire _al_u1622_o;
  wire _al_u1623_o;
  wire _al_u1624_o;
  wire _al_u1625_o;
  wire _al_u1626_o;
  wire _al_u1627_o;
  wire _al_u1628_o;
  wire _al_u1629_o;
  wire _al_u1630_o;
  wire _al_u1631_o;
  wire _al_u1632_o;
  wire _al_u1633_o;
  wire _al_u1634_o;
  wire _al_u1635_o;
  wire _al_u1636_o;
  wire _al_u1638_o;
  wire _al_u1639_o;
  wire _al_u1640_o;
  wire _al_u1641_o;
  wire _al_u1642_o;
  wire _al_u1643_o;
  wire _al_u1644_o;
  wire _al_u1645_o;
  wire _al_u1646_o;
  wire _al_u1647_o;
  wire _al_u1648_o;
  wire _al_u1649_o;
  wire _al_u1650_o;
  wire _al_u1651_o;
  wire _al_u1652_o;
  wire _al_u1653_o;
  wire _al_u1654_o;
  wire _al_u1655_o;
  wire _al_u1656_o;
  wire _al_u1657_o;
  wire _al_u1659_o;
  wire _al_u1660_o;
  wire _al_u1661_o;
  wire _al_u1662_o;
  wire _al_u1663_o;
  wire _al_u1664_o;
  wire _al_u1665_o;
  wire _al_u1666_o;
  wire _al_u1667_o;
  wire _al_u1668_o;
  wire _al_u1669_o;
  wire _al_u1670_o;
  wire _al_u1671_o;
  wire _al_u1672_o;
  wire _al_u1673_o;
  wire _al_u1674_o;
  wire _al_u1675_o;
  wire _al_u1676_o;
  wire _al_u1677_o;
  wire _al_u1678_o;
  wire _al_u1680_o;
  wire _al_u1681_o;
  wire _al_u1682_o;
  wire _al_u1683_o;
  wire _al_u1684_o;
  wire _al_u1685_o;
  wire _al_u1686_o;
  wire _al_u1687_o;
  wire _al_u1688_o;
  wire _al_u1689_o;
  wire _al_u1690_o;
  wire _al_u1691_o;
  wire _al_u1692_o;
  wire _al_u1693_o;
  wire _al_u1694_o;
  wire _al_u1695_o;
  wire _al_u1696_o;
  wire _al_u1697_o;
  wire _al_u1698_o;
  wire _al_u1699_o;
  wire _al_u1701_o;
  wire _al_u1702_o;
  wire _al_u1703_o;
  wire _al_u1704_o;
  wire _al_u1705_o;
  wire _al_u1706_o;
  wire _al_u1707_o;
  wire _al_u1708_o;
  wire _al_u1709_o;
  wire _al_u1710_o;
  wire _al_u1711_o;
  wire _al_u1712_o;
  wire _al_u1713_o;
  wire _al_u1714_o;
  wire _al_u1715_o;
  wire _al_u1716_o;
  wire _al_u1717_o;
  wire _al_u1718_o;
  wire _al_u1719_o;
  wire _al_u1720_o;
  wire _al_u1722_o;
  wire _al_u1723_o;
  wire _al_u1724_o;
  wire _al_u1725_o;
  wire _al_u1727_o;
  wire _al_u1728_o;
  wire _al_u1729_o;
  wire _al_u1730_o;
  wire _al_u1733_o;
  wire _al_u1734_o;
  wire _al_u1735_o;
  wire _al_u1736_o;
  wire _al_u1737_o;
  wire _al_u1739_o;
  wire _al_u1740_o;
  wire _al_u1742_o;
  wire _al_u1743_o;
  wire _al_u1744_o;
  wire _al_u1745_o;
  wire _al_u1747_o;
  wire _al_u1783_o;
  wire _al_u1784_o;
  wire _al_u1785_o;
  wire _al_u1786_o;
  wire _al_u1788_o;
  wire _al_u1789_o;
  wire _al_u1790_o;
  wire _al_u1791_o;
  wire _al_u1792_o;
  wire _al_u1793_o;
  wire _al_u1796_o;
  wire _al_u1797_o;
  wire _al_u1798_o;
  wire _al_u1800_o;
  wire _al_u1801_o;
  wire _al_u1802_o;
  wire _al_u1803_o;
  wire _al_u1806_o;
  wire _al_u1808_o;
  wire _al_u1811_o;
  wire _al_u1814_o;
  wire _al_u1817_o;
  wire _al_u1820_o;
  wire _al_u1823_o;
  wire _al_u1826_o;
  wire _al_u1829_o;
  wire _al_u1832_o;
  wire _al_u1835_o;
  wire _al_u1838_o;
  wire _al_u1841_o;
  wire _al_u1844_o;
  wire _al_u1847_o;
  wire _al_u1850_o;
  wire _al_u1853_o;
  wire _al_u1856_o;
  wire _al_u1859_o;
  wire _al_u1862_o;
  wire _al_u1865_o;
  wire _al_u1868_o;
  wire _al_u1871_o;
  wire _al_u1874_o;
  wire _al_u1877_o;
  wire _al_u1880_o;
  wire _al_u1883_o;
  wire _al_u1886_o;
  wire _al_u1889_o;
  wire _al_u1892_o;
  wire _al_u1895_o;
  wire _al_u1898_o;
  wire _al_u1902_o;
  wire _al_u1903_o;
  wire _al_u1904_o;
  wire _al_u1906_o;
  wire _al_u1908_o;
  wire _al_u1916_o;
  wire _al_u1917_o;
  wire _al_u1918_o;
  wire _al_u1935_o;
  wire _al_u1940_o;
  wire _al_u1944_o;
  wire _al_u1947_o;
  wire _al_u1948_o;
  wire _al_u1950_o;
  wire _al_u1956_o;
  wire _al_u1958_o;
  wire _al_u1960_o;
  wire _al_u1962_o;
  wire _al_u1965_o;
  wire _al_u1967_o;
  wire _al_u1968_o;
  wire _al_u1969_o;
  wire _al_u1970_o;
  wire _al_u1973_o;
  wire _al_u1974_o;
  wire _al_u1975_o;
  wire _al_u1976_o;
  wire _al_u1979_o;
  wire _al_u1983_o;
  wire _al_u1984_o;
  wire _al_u1985_o;
  wire _al_u1987_o;
  wire _al_u1990_o;
  wire _al_u1993_o;
  wire _al_u1996_o;
  wire _al_u1999_o;
  wire _al_u2000_o;
  wire _al_u2002_o;
  wire _al_u2005_o;
  wire _al_u2007_o;
  wire _al_u2009_o;
  wire _al_u2010_o;
  wire _al_u2012_o;
  wire _al_u2015_o;
  wire _al_u2018_o;
  wire _al_u2021_o;
  wire _al_u2024_o;
  wire _al_u2027_o;
  wire _al_u2030_o;
  wire _al_u2033_o;
  wire _al_u2036_o;
  wire _al_u2039_o;
  wire _al_u2042_o;
  wire _al_u2045_o;
  wire _al_u2048_o;
  wire _al_u2051_o;
  wire _al_u2054_o;
  wire _al_u2057_o;
  wire _al_u2060_o;
  wire _al_u2063_o;
  wire _al_u2066_o;
  wire _al_u2069_o;
  wire _al_u2072_o;
  wire _al_u2073_o;
  wire _al_u2075_o;
  wire _al_u2076_o;
  wire _al_u2078_o;
  wire _al_u2080_o;
  wire _al_u2092_o;
  wire _al_u2093_o;
  wire _al_u2095_o;
  wire _al_u2096_o;
  wire _al_u2097_o;
  wire _al_u2098_o;
  wire _al_u2099_o;
  wire _al_u2100_o;
  wire _al_u2101_o;
  wire _al_u2102_o;
  wire _al_u2103_o;
  wire _al_u2104_o;
  wire _al_u2105_o;
  wire _al_u2106_o;
  wire _al_u2107_o;
  wire _al_u2109_o;
  wire _al_u2111_o;
  wire _al_u2113_o;
  wire _al_u2115_o;
  wire _al_u2117_o;
  wire _al_u2119_o;
  wire _al_u2124_o;
  wire _al_u2126_o;
  wire _al_u2128_o;
  wire _al_u2130_o;
  wire _al_u2133_o;
  wire _al_u2136_o;
  wire _al_u2137_o;
  wire _al_u2140_o;
  wire _al_u2143_o;
  wire _al_u2144_o;
  wire _al_u2145_o;
  wire _al_u2146_o;
  wire _al_u2147_o;
  wire _al_u2150_o;
  wire _al_u2153_o;
  wire _al_u2154_o;
  wire _al_u2157_o;
  wire _al_u2159_o;
  wire _al_u2161_o;
  wire _al_u2162_o;
  wire _al_u2163_o;
  wire _al_u2165_o;
  wire _al_u2166_o;
  wire _al_u2168_o;
  wire _al_u2169_o;
  wire _al_u2170_o;
  wire _al_u2172_o;
  wire _al_u2175_o;
  wire _al_u2178_o;
  wire _al_u2179_o;
  wire _al_u2182_o;
  wire _al_u2184_o;
  wire _al_u2185_o;
  wire _al_u2186_o;
  wire _al_u2187_o;
  wire _al_u2188_o;
  wire _al_u2191_o;
  wire _al_u2194_o;
  wire _al_u2195_o;
  wire _al_u2198_o;
  wire _al_u2201_o;
  wire _al_u2202_o;
  wire _al_u2203_o;
  wire _al_u2208_o;
  wire _al_u2209_o;
  wire _al_u2210_o;
  wire _al_u2212_o;
  wire _al_u2213_o;
  wire _al_u2214_o;
  wire _al_u2215_o;
  wire _al_u2216_o;
  wire _al_u2218_o;
  wire _al_u2219_o;
  wire _al_u2220_o;
  wire _al_u2221_o;
  wire _al_u2222_o;
  wire _al_u2223_o;
  wire _al_u2224_o;
  wire _al_u2225_o;
  wire _al_u2226_o;
  wire _al_u2227_o;
  wire _al_u2229_o;
  wire _al_u2232_o;
  wire _al_u2233_o;
  wire _al_u2234_o;
  wire _al_u2236_o;
  wire _al_u2237_o;
  wire _al_u2238_o;
  wire _al_u2239_o;
  wire _al_u2240_o;
  wire _al_u2241_o;
  wire _al_u2242_o;
  wire _al_u2243_o;
  wire _al_u2244_o;
  wire _al_u2245_o;
  wire _al_u2246_o;
  wire _al_u2247_o;
  wire _al_u2248_o;
  wire _al_u2249_o;
  wire _al_u2250_o;
  wire _al_u2252_o;
  wire _al_u2255_o;
  wire _al_u2256_o;
  wire _al_u2257_o;
  wire _al_u2259_o;
  wire _al_u2260_o;
  wire _al_u2262_o;
  wire _al_u2263_o;
  wire _al_u2264_o;
  wire _al_u2265_o;
  wire _al_u2266_o;
  wire _al_u2267_o;
  wire _al_u2269_o;
  wire _al_u2270_o;
  wire _al_u2272_o;
  wire _al_u2273_o;
  wire _al_u2274_o;
  wire _al_u2276_o;
  wire _al_u2277_o;
  wire _al_u2279_o;
  wire _al_u2280_o;
  wire _al_u2281_o;
  wire _al_u2282_o;
  wire _al_u2283_o;
  wire _al_u2284_o;
  wire _al_u2286_o;
  wire _al_u2287_o;
  wire _al_u2289_o;
  wire _al_u2290_o;
  wire _al_u2291_o;
  wire _al_u2293_o;
  wire _al_u2294_o;
  wire _al_u2296_o;
  wire _al_u2297_o;
  wire _al_u2298_o;
  wire _al_u2299_o;
  wire _al_u2300_o;
  wire _al_u2301_o;
  wire _al_u2303_o;
  wire _al_u2304_o;
  wire _al_u2306_o;
  wire _al_u2307_o;
  wire _al_u2308_o;
  wire _al_u2310_o;
  wire _al_u2311_o;
  wire _al_u2312_o;
  wire _al_u2313_o;
  wire _al_u2314_o;
  wire _al_u2315_o;
  wire _al_u2316_o;
  wire _al_u2317_o;
  wire _al_u2319_o;
  wire _al_u2320_o;
  wire _al_u2322_o;
  wire _al_u2323_o;
  wire _al_u2324_o;
  wire _al_u2327_o;
  wire _al_u2328_o;
  wire _al_u2329_o;
  wire _al_u2330_o;
  wire _al_u2332_o;
  wire _al_u2333_o;
  wire _al_u2334_o;
  wire _al_u2335_o;
  wire _al_u2336_o;
  wire _al_u2337_o;
  wire _al_u2340_o;
  wire _al_u2341_o;
  wire _al_u2342_o;
  wire _al_u2343_o;
  wire _al_u2345_o;
  wire _al_u2346_o;
  wire _al_u2347_o;
  wire _al_u2348_o;
  wire _al_u2349_o;
  wire _al_u2350_o;
  wire _al_u2353_o;
  wire _al_u2354_o;
  wire _al_u2355_o;
  wire _al_u2356_o;
  wire _al_u2358_o;
  wire _al_u2359_o;
  wire _al_u2360_o;
  wire _al_u2361_o;
  wire _al_u2362_o;
  wire _al_u2363_o;
  wire _al_u2366_o;
  wire _al_u2367_o;
  wire _al_u2368_o;
  wire _al_u2369_o;
  wire _al_u2371_o;
  wire _al_u2372_o;
  wire _al_u2373_o;
  wire _al_u2374_o;
  wire _al_u2375_o;
  wire _al_u2376_o;
  wire _al_u2378_o;
  wire _al_u2380_o;
  wire _al_u2381_o;
  wire _al_u2383_o;
  wire _al_u2384_o;
  wire _al_u2385_o;
  wire _al_u2386_o;
  wire _al_u2387_o;
  wire _al_u2388_o;
  wire _al_u2390_o;
  wire _al_u2392_o;
  wire _al_u2393_o;
  wire _al_u2395_o;
  wire _al_u2396_o;
  wire _al_u2397_o;
  wire _al_u2398_o;
  wire _al_u2399_o;
  wire _al_u2400_o;
  wire _al_u2403_o;
  wire _al_u2404_o;
  wire _al_u2405_o;
  wire _al_u2406_o;
  wire _al_u2408_o;
  wire _al_u2409_o;
  wire _al_u2410_o;
  wire _al_u2411_o;
  wire _al_u2412_o;
  wire _al_u2413_o;
  wire _al_u2415_o;
  wire _al_u2416_o;
  wire _al_u2417_o;
  wire _al_u2418_o;
  wire _al_u2420_o;
  wire _al_u2421_o;
  wire _al_u2422_o;
  wire _al_u2423_o;
  wire _al_u2424_o;
  wire _al_u2425_o;
  wire _al_u2427_o;
  wire _al_u2429_o;
  wire _al_u2430_o;
  wire _al_u2431_o;
  wire _al_u2432_o;
  wire _al_u2433_o;
  wire _al_u2434_o;
  wire _al_u2435_o;
  wire _al_u2436_o;
  wire _al_u2438_o;
  wire _al_u2439_o;
  wire _al_u2440_o;
  wire _al_u2442_o;
  wire _al_u2443_o;
  wire _al_u2444_o;
  wire _al_u2445_o;
  wire _al_u2446_o;
  wire _al_u2448_o;
  wire _al_u2449_o;
  wire _al_u2450_o;
  wire _al_u2452_o;
  wire _al_u2453_o;
  wire _al_u2454_o;
  wire _al_u2455_o;
  wire _al_u2456_o;
  wire _al_u2458_o;
  wire _al_u2459_o;
  wire _al_u2460_o;
  wire _al_u2462_o;
  wire _al_u2463_o;
  wire _al_u2464_o;
  wire _al_u2465_o;
  wire _al_u2466_o;
  wire _al_u2468_o;
  wire _al_u2469_o;
  wire _al_u2470_o;
  wire _al_u2472_o;
  wire _al_u2473_o;
  wire _al_u2474_o;
  wire _al_u2475_o;
  wire _al_u2476_o;
  wire _al_u2478_o;
  wire _al_u2479_o;
  wire _al_u2480_o;
  wire _al_u2482_o;
  wire _al_u2483_o;
  wire _al_u2484_o;
  wire _al_u2485_o;
  wire _al_u2486_o;
  wire _al_u2488_o;
  wire _al_u2489_o;
  wire _al_u2490_o;
  wire _al_u2492_o;
  wire _al_u2493_o;
  wire _al_u2494_o;
  wire _al_u2495_o;
  wire _al_u2496_o;
  wire _al_u2498_o;
  wire _al_u2499_o;
  wire _al_u2500_o;
  wire _al_u2502_o;
  wire _al_u2503_o;
  wire _al_u2504_o;
  wire _al_u2505_o;
  wire _al_u2506_o;
  wire _al_u2508_o;
  wire _al_u2509_o;
  wire _al_u2510_o;
  wire _al_u2512_o;
  wire _al_u2513_o;
  wire _al_u2514_o;
  wire _al_u2515_o;
  wire _al_u2516_o;
  wire _al_u251_o;
  wire _al_u2520_o;
  wire _al_u2521_o;
  wire _al_u2522_o;
  wire _al_u2523_o;
  wire _al_u2524_o;
  wire _al_u2525_o;
  wire _al_u2526_o;
  wire _al_u252_o;
  wire _al_u2530_o;
  wire _al_u2531_o;
  wire _al_u2532_o;
  wire _al_u2533_o;
  wire _al_u2534_o;
  wire _al_u2535_o;
  wire _al_u2536_o;
  wire _al_u2538_o;
  wire _al_u2539_o;
  wire _al_u2540_o;
  wire _al_u2541_o;
  wire _al_u2543_o;
  wire _al_u2544_o;
  wire _al_u2545_o;
  wire _al_u2546_o;
  wire _al_u2547_o;
  wire _al_u254_o;
  wire _al_u2551_o;
  wire _al_u2552_o;
  wire _al_u2553_o;
  wire _al_u2554_o;
  wire _al_u2555_o;
  wire _al_u2556_o;
  wire _al_u2560_o;
  wire _al_u2561_o;
  wire _al_u2562_o;
  wire _al_u2563_o;
  wire _al_u2564_o;
  wire _al_u2565_o;
  wire _al_u2567_o;
  wire _al_u2568_o;
  wire _al_u2569_o;
  wire _al_u256_o;
  wire _al_u2570_o;
  wire _al_u2571_o;
  wire _al_u2572_o;
  wire _al_u2573_o;
  wire _al_u2574_o;
  wire _al_u2575_o;
  wire _al_u2576_o;
  wire _al_u2577_o;
  wire _al_u2580_o;
  wire _al_u2581_o;
  wire _al_u2582_o;
  wire _al_u2583_o;
  wire _al_u2584_o;
  wire _al_u2585_o;
  wire _al_u2586_o;
  wire _al_u2587_o;
  wire _al_u2589_o;
  wire _al_u2590_o;
  wire _al_u2591_o;
  wire _al_u2592_o;
  wire _al_u2593_o;
  wire _al_u2594_o;
  wire _al_u2595_o;
  wire _al_u2596_o;
  wire _al_u2597_o;
  wire _al_u2598_o;
  wire _al_u2599_o;
  wire _al_u2600_o;
  wire _al_u2601_o;
  wire _al_u2602_o;
  wire _al_u2604_o;
  wire _al_u2606_o;
  wire _al_u2607_o;
  wire _al_u2608_o;
  wire _al_u2609_o;
  wire _al_u2610_o;
  wire _al_u2611_o;
  wire _al_u2613_o;
  wire _al_u2614_o;
  wire _al_u2615_o;
  wire _al_u2616_o;
  wire _al_u2617_o;
  wire _al_u2619_o;
  wire _al_u2621_o;
  wire _al_u2623_o;
  wire _al_u2625_o;
  wire _al_u2627_o;
  wire _al_u2629_o;
  wire _al_u2631_o;
  wire _al_u2633_o;
  wire _al_u2635_o;
  wire _al_u2637_o;
  wire _al_u2639_o;
  wire _al_u2641_o;
  wire _al_u2643_o;
  wire _al_u2645_o;
  wire _al_u2647_o;
  wire _al_u2649_o;
  wire _al_u2651_o;
  wire _al_u2653_o;
  wire _al_u2655_o;
  wire _al_u2657_o;
  wire _al_u2659_o;
  wire _al_u2661_o;
  wire _al_u2663_o;
  wire _al_u2665_o;
  wire _al_u2667_o;
  wire _al_u2669_o;
  wire _al_u2671_o;
  wire _al_u2673_o;
  wire _al_u2675_o;
  wire _al_u2677_o;
  wire _al_u2679_o;
  wire _al_u2680_o;
  wire _al_u2681_o;
  wire _al_u2683_o;
  wire _al_u2684_o;
  wire _al_u2686_o;
  wire _al_u2687_o;
  wire _al_u2688_o;
  wire _al_u2689_o;
  wire _al_u2690_o;
  wire _al_u2692_o;
  wire _al_u2693_o;
  wire _al_u2695_o;
  wire _al_u2697_o;
  wire _al_u2699_o;
  wire _al_u2701_o;
  wire _al_u2703_o;
  wire _al_u2705_o;
  wire _al_u2707_o;
  wire _al_u2708_o;
  wire _al_u2709_o;
  wire _al_u2710_o;
  wire _al_u2711_o;
  wire _al_u2713_o;
  wire _al_u2714_o;
  wire _al_u2716_o;
  wire _al_u2718_o;
  wire _al_u2720_o;
  wire _al_u2722_o;
  wire _al_u2724_o;
  wire _al_u2726_o;
  wire _al_u2728_o;
  wire _al_u2729_o;
  wire _al_u2730_o;
  wire _al_u2732_o;
  wire _al_u2733_o;
  wire _al_u2735_o;
  wire _al_u2736_o;
  wire _al_u2737_o;
  wire _al_u2739_o;
  wire _al_u2740_o;
  wire _al_u2742_o;
  wire _al_u2744_o;
  wire _al_u2745_o;
  wire _al_u2747_o;
  wire _al_u2748_o;
  wire _al_u2749_o;
  wire _al_u2751_o;
  wire _al_u2752_o;
  wire _al_u2754_o;
  wire _al_u2756_o;
  wire _al_u2758_o;
  wire _al_u2760_o;
  wire _al_u2762_o;
  wire _al_u2764_o;
  wire _al_u2766_o;
  wire _al_u2767_o;
  wire _al_u2768_o;
  wire _al_u2769_o;
  wire _al_u2770_o;
  wire _al_u2771_o;
  wire _al_u2772_o;
  wire _al_u2773_o;
  wire _al_u2774_o;
  wire _al_u2775_o;
  wire _al_u2776_o;
  wire _al_u2777_o;
  wire _al_u2778_o;
  wire _al_u2779_o;
  wire _al_u2780_o;
  wire _al_u2781_o;
  wire _al_u2782_o;
  wire _al_u2783_o;
  wire _al_u2784_o;
  wire _al_u2785_o;
  wire _al_u2786_o;
  wire _al_u2787_o;
  wire _al_u2788_o;
  wire _al_u2789_o;
  wire _al_u2790_o;
  wire _al_u2791_o;
  wire _al_u2792_o;
  wire _al_u2793_o;
  wire _al_u2794_o;
  wire _al_u2795_o;
  wire _al_u2796_o;
  wire _al_u2798_o;
  wire _al_u2799_o;
  wire _al_u2800_o;
  wire _al_u2801_o;
  wire _al_u2802_o;
  wire _al_u2803_o;
  wire _al_u2806_o;
  wire _al_u2807_o;
  wire _al_u2808_o;
  wire _al_u2810_o;
  wire _al_u2811_o;
  wire _al_u2812_o;
  wire _al_u2814_o;
  wire _al_u2815_o;
  wire _al_u2817_o;
  wire _al_u2819_o;
  wire _al_u2821_o;
  wire _al_u2822_o;
  wire _al_u2824_o;
  wire _al_u2826_o;
  wire _al_u2828_o;
  wire _al_u2829_o;
  wire _al_u2831_o;
  wire _al_u2833_o;
  wire _al_u2834_o;
  wire _al_u2836_o;
  wire _al_u2838_o;
  wire _al_u2840_o;
  wire _al_u2841_o;
  wire _al_u2843_o;
  wire _al_u2844_o;
  wire _al_u2846_o;
  wire _al_u2847_o;
  wire _al_u2849_o;
  wire _al_u2850_o;
  wire _al_u2852_o;
  wire _al_u2854_o;
  wire _al_u2856_o;
  wire _al_u2857_o;
  wire _al_u2859_o;
  wire _al_u2860_o;
  wire _al_u2862_o;
  wire _al_u2864_o;
  wire _al_u2866_o;
  wire _al_u2868_o;
  wire _al_u2869_o;
  wire _al_u2871_o;
  wire _al_u2872_o;
  wire _al_u2874_o;
  wire _al_u2875_o;
  wire _al_u2877_o;
  wire _al_u2878_o;
  wire _al_u2880_o;
  wire _al_u2882_o;
  wire _al_u2883_o;
  wire _al_u2885_o;
  wire _al_u2887_o;
  wire _al_u2888_o;
  wire _al_u2890_o;
  wire _al_u290_o;
  wire _al_u328_o;
  wire _al_u329_o;
  wire _al_u330_o;
  wire _al_u331_o;
  wire _al_u333_o;
  wire _al_u334_o;
  wire _al_u335_o;
  wire _al_u336_o;
  wire _al_u337_o;
  wire _al_u338_o;
  wire _al_u339_o;
  wire _al_u340_o;
  wire _al_u341_o;
  wire _al_u342_o;
  wire _al_u343_o;
  wire _al_u344_o;
  wire _al_u345_o;
  wire _al_u346_o;
  wire _al_u347_o;
  wire _al_u348_o;
  wire _al_u349_o;
  wire _al_u350_o;
  wire _al_u351_o;
  wire _al_u352_o;
  wire _al_u353_o;
  wire _al_u355_o;
  wire _al_u356_o;
  wire _al_u357_o;
  wire _al_u358_o;
  wire _al_u359_o;
  wire _al_u360_o;
  wire _al_u361_o;
  wire _al_u362_o;
  wire _al_u363_o;
  wire _al_u364_o;
  wire _al_u365_o;
  wire _al_u366_o;
  wire _al_u367_o;
  wire _al_u368_o;
  wire _al_u369_o;
  wire _al_u370_o;
  wire _al_u371_o;
  wire _al_u372_o;
  wire _al_u373_o;
  wire _al_u374_o;
  wire _al_u376_o;
  wire _al_u377_o;
  wire _al_u378_o;
  wire _al_u379_o;
  wire _al_u380_o;
  wire _al_u381_o;
  wire _al_u382_o;
  wire _al_u383_o;
  wire _al_u384_o;
  wire _al_u385_o;
  wire _al_u386_o;
  wire _al_u387_o;
  wire _al_u388_o;
  wire _al_u389_o;
  wire _al_u390_o;
  wire _al_u391_o;
  wire _al_u392_o;
  wire _al_u393_o;
  wire _al_u394_o;
  wire _al_u395_o;
  wire _al_u397_o;
  wire _al_u398_o;
  wire _al_u399_o;
  wire _al_u400_o;
  wire _al_u401_o;
  wire _al_u402_o;
  wire _al_u403_o;
  wire _al_u404_o;
  wire _al_u405_o;
  wire _al_u406_o;
  wire _al_u407_o;
  wire _al_u408_o;
  wire _al_u409_o;
  wire _al_u410_o;
  wire _al_u411_o;
  wire _al_u412_o;
  wire _al_u413_o;
  wire _al_u414_o;
  wire _al_u415_o;
  wire _al_u416_o;
  wire _al_u418_o;
  wire _al_u419_o;
  wire _al_u420_o;
  wire _al_u421_o;
  wire _al_u422_o;
  wire _al_u423_o;
  wire _al_u424_o;
  wire _al_u425_o;
  wire _al_u426_o;
  wire _al_u427_o;
  wire _al_u428_o;
  wire _al_u429_o;
  wire _al_u430_o;
  wire _al_u431_o;
  wire _al_u432_o;
  wire _al_u433_o;
  wire _al_u434_o;
  wire _al_u435_o;
  wire _al_u436_o;
  wire _al_u437_o;
  wire _al_u439_o;
  wire _al_u440_o;
  wire _al_u441_o;
  wire _al_u442_o;
  wire _al_u443_o;
  wire _al_u444_o;
  wire _al_u445_o;
  wire _al_u446_o;
  wire _al_u447_o;
  wire _al_u448_o;
  wire _al_u449_o;
  wire _al_u450_o;
  wire _al_u451_o;
  wire _al_u452_o;
  wire _al_u453_o;
  wire _al_u454_o;
  wire _al_u455_o;
  wire _al_u456_o;
  wire _al_u457_o;
  wire _al_u458_o;
  wire _al_u460_o;
  wire _al_u461_o;
  wire _al_u462_o;
  wire _al_u463_o;
  wire _al_u464_o;
  wire _al_u465_o;
  wire _al_u466_o;
  wire _al_u467_o;
  wire _al_u468_o;
  wire _al_u469_o;
  wire _al_u470_o;
  wire _al_u471_o;
  wire _al_u472_o;
  wire _al_u473_o;
  wire _al_u474_o;
  wire _al_u475_o;
  wire _al_u476_o;
  wire _al_u477_o;
  wire _al_u478_o;
  wire _al_u479_o;
  wire _al_u481_o;
  wire _al_u482_o;
  wire _al_u483_o;
  wire _al_u484_o;
  wire _al_u485_o;
  wire _al_u486_o;
  wire _al_u487_o;
  wire _al_u488_o;
  wire _al_u489_o;
  wire _al_u490_o;
  wire _al_u491_o;
  wire _al_u492_o;
  wire _al_u493_o;
  wire _al_u494_o;
  wire _al_u495_o;
  wire _al_u496_o;
  wire _al_u497_o;
  wire _al_u498_o;
  wire _al_u499_o;
  wire _al_u500_o;
  wire _al_u502_o;
  wire _al_u503_o;
  wire _al_u504_o;
  wire _al_u505_o;
  wire _al_u506_o;
  wire _al_u507_o;
  wire _al_u508_o;
  wire _al_u509_o;
  wire _al_u510_o;
  wire _al_u511_o;
  wire _al_u512_o;
  wire _al_u513_o;
  wire _al_u514_o;
  wire _al_u515_o;
  wire _al_u516_o;
  wire _al_u517_o;
  wire _al_u518_o;
  wire _al_u519_o;
  wire _al_u520_o;
  wire _al_u521_o;
  wire _al_u523_o;
  wire _al_u524_o;
  wire _al_u525_o;
  wire _al_u526_o;
  wire _al_u527_o;
  wire _al_u528_o;
  wire _al_u529_o;
  wire _al_u530_o;
  wire _al_u531_o;
  wire _al_u532_o;
  wire _al_u533_o;
  wire _al_u534_o;
  wire _al_u535_o;
  wire _al_u536_o;
  wire _al_u537_o;
  wire _al_u538_o;
  wire _al_u539_o;
  wire _al_u540_o;
  wire _al_u541_o;
  wire _al_u542_o;
  wire _al_u544_o;
  wire _al_u545_o;
  wire _al_u546_o;
  wire _al_u547_o;
  wire _al_u548_o;
  wire _al_u549_o;
  wire _al_u550_o;
  wire _al_u551_o;
  wire _al_u552_o;
  wire _al_u553_o;
  wire _al_u554_o;
  wire _al_u555_o;
  wire _al_u556_o;
  wire _al_u557_o;
  wire _al_u558_o;
  wire _al_u559_o;
  wire _al_u560_o;
  wire _al_u561_o;
  wire _al_u562_o;
  wire _al_u563_o;
  wire _al_u565_o;
  wire _al_u566_o;
  wire _al_u567_o;
  wire _al_u568_o;
  wire _al_u569_o;
  wire _al_u570_o;
  wire _al_u571_o;
  wire _al_u572_o;
  wire _al_u573_o;
  wire _al_u574_o;
  wire _al_u575_o;
  wire _al_u576_o;
  wire _al_u577_o;
  wire _al_u578_o;
  wire _al_u579_o;
  wire _al_u580_o;
  wire _al_u581_o;
  wire _al_u582_o;
  wire _al_u583_o;
  wire _al_u584_o;
  wire _al_u586_o;
  wire _al_u587_o;
  wire _al_u588_o;
  wire _al_u589_o;
  wire _al_u590_o;
  wire _al_u591_o;
  wire _al_u592_o;
  wire _al_u593_o;
  wire _al_u594_o;
  wire _al_u595_o;
  wire _al_u596_o;
  wire _al_u597_o;
  wire _al_u598_o;
  wire _al_u599_o;
  wire _al_u600_o;
  wire _al_u601_o;
  wire _al_u602_o;
  wire _al_u603_o;
  wire _al_u604_o;
  wire _al_u605_o;
  wire _al_u607_o;
  wire _al_u608_o;
  wire _al_u609_o;
  wire _al_u610_o;
  wire _al_u611_o;
  wire _al_u612_o;
  wire _al_u613_o;
  wire _al_u614_o;
  wire _al_u615_o;
  wire _al_u616_o;
  wire _al_u617_o;
  wire _al_u618_o;
  wire _al_u619_o;
  wire _al_u620_o;
  wire _al_u621_o;
  wire _al_u622_o;
  wire _al_u623_o;
  wire _al_u624_o;
  wire _al_u625_o;
  wire _al_u626_o;
  wire _al_u628_o;
  wire _al_u629_o;
  wire _al_u630_o;
  wire _al_u631_o;
  wire _al_u632_o;
  wire _al_u633_o;
  wire _al_u634_o;
  wire _al_u635_o;
  wire _al_u636_o;
  wire _al_u637_o;
  wire _al_u638_o;
  wire _al_u639_o;
  wire _al_u640_o;
  wire _al_u641_o;
  wire _al_u642_o;
  wire _al_u643_o;
  wire _al_u644_o;
  wire _al_u645_o;
  wire _al_u646_o;
  wire _al_u647_o;
  wire _al_u649_o;
  wire _al_u650_o;
  wire _al_u651_o;
  wire _al_u652_o;
  wire _al_u653_o;
  wire _al_u654_o;
  wire _al_u655_o;
  wire _al_u656_o;
  wire _al_u657_o;
  wire _al_u658_o;
  wire _al_u659_o;
  wire _al_u660_o;
  wire _al_u661_o;
  wire _al_u662_o;
  wire _al_u663_o;
  wire _al_u664_o;
  wire _al_u665_o;
  wire _al_u666_o;
  wire _al_u667_o;
  wire _al_u668_o;
  wire _al_u670_o;
  wire _al_u671_o;
  wire _al_u672_o;
  wire _al_u673_o;
  wire _al_u674_o;
  wire _al_u675_o;
  wire _al_u676_o;
  wire _al_u677_o;
  wire _al_u678_o;
  wire _al_u679_o;
  wire _al_u680_o;
  wire _al_u681_o;
  wire _al_u682_o;
  wire _al_u683_o;
  wire _al_u684_o;
  wire _al_u685_o;
  wire _al_u686_o;
  wire _al_u687_o;
  wire _al_u688_o;
  wire _al_u689_o;
  wire _al_u691_o;
  wire _al_u692_o;
  wire _al_u693_o;
  wire _al_u694_o;
  wire _al_u695_o;
  wire _al_u696_o;
  wire _al_u697_o;
  wire _al_u698_o;
  wire _al_u699_o;
  wire _al_u700_o;
  wire _al_u701_o;
  wire _al_u702_o;
  wire _al_u703_o;
  wire _al_u704_o;
  wire _al_u705_o;
  wire _al_u706_o;
  wire _al_u707_o;
  wire _al_u708_o;
  wire _al_u709_o;
  wire _al_u710_o;
  wire _al_u712_o;
  wire _al_u713_o;
  wire _al_u714_o;
  wire _al_u715_o;
  wire _al_u716_o;
  wire _al_u717_o;
  wire _al_u718_o;
  wire _al_u719_o;
  wire _al_u720_o;
  wire _al_u721_o;
  wire _al_u722_o;
  wire _al_u723_o;
  wire _al_u724_o;
  wire _al_u725_o;
  wire _al_u726_o;
  wire _al_u727_o;
  wire _al_u728_o;
  wire _al_u729_o;
  wire _al_u730_o;
  wire _al_u731_o;
  wire _al_u733_o;
  wire _al_u734_o;
  wire _al_u735_o;
  wire _al_u736_o;
  wire _al_u737_o;
  wire _al_u738_o;
  wire _al_u739_o;
  wire _al_u740_o;
  wire _al_u741_o;
  wire _al_u742_o;
  wire _al_u743_o;
  wire _al_u744_o;
  wire _al_u745_o;
  wire _al_u746_o;
  wire _al_u747_o;
  wire _al_u748_o;
  wire _al_u749_o;
  wire _al_u750_o;
  wire _al_u751_o;
  wire _al_u752_o;
  wire _al_u754_o;
  wire _al_u755_o;
  wire _al_u756_o;
  wire _al_u757_o;
  wire _al_u758_o;
  wire _al_u759_o;
  wire _al_u760_o;
  wire _al_u761_o;
  wire _al_u762_o;
  wire _al_u763_o;
  wire _al_u764_o;
  wire _al_u765_o;
  wire _al_u766_o;
  wire _al_u767_o;
  wire _al_u768_o;
  wire _al_u769_o;
  wire _al_u770_o;
  wire _al_u771_o;
  wire _al_u772_o;
  wire _al_u773_o;
  wire _al_u775_o;
  wire _al_u776_o;
  wire _al_u777_o;
  wire _al_u778_o;
  wire _al_u779_o;
  wire _al_u780_o;
  wire _al_u781_o;
  wire _al_u782_o;
  wire _al_u783_o;
  wire _al_u784_o;
  wire _al_u785_o;
  wire _al_u786_o;
  wire _al_u787_o;
  wire _al_u788_o;
  wire _al_u789_o;
  wire _al_u790_o;
  wire _al_u791_o;
  wire _al_u792_o;
  wire _al_u793_o;
  wire _al_u794_o;
  wire _al_u796_o;
  wire _al_u797_o;
  wire _al_u798_o;
  wire _al_u799_o;
  wire _al_u800_o;
  wire _al_u801_o;
  wire _al_u802_o;
  wire _al_u803_o;
  wire _al_u804_o;
  wire _al_u805_o;
  wire _al_u806_o;
  wire _al_u807_o;
  wire _al_u808_o;
  wire _al_u809_o;
  wire _al_u810_o;
  wire _al_u811_o;
  wire _al_u812_o;
  wire _al_u813_o;
  wire _al_u814_o;
  wire _al_u815_o;
  wire _al_u817_o;
  wire _al_u818_o;
  wire _al_u819_o;
  wire _al_u820_o;
  wire _al_u821_o;
  wire _al_u822_o;
  wire _al_u823_o;
  wire _al_u824_o;
  wire _al_u825_o;
  wire _al_u826_o;
  wire _al_u827_o;
  wire _al_u828_o;
  wire _al_u829_o;
  wire _al_u830_o;
  wire _al_u831_o;
  wire _al_u832_o;
  wire _al_u833_o;
  wire _al_u834_o;
  wire _al_u835_o;
  wire _al_u836_o;
  wire _al_u838_o;
  wire _al_u839_o;
  wire _al_u840_o;
  wire _al_u841_o;
  wire _al_u842_o;
  wire _al_u843_o;
  wire _al_u844_o;
  wire _al_u845_o;
  wire _al_u846_o;
  wire _al_u847_o;
  wire _al_u848_o;
  wire _al_u849_o;
  wire _al_u850_o;
  wire _al_u851_o;
  wire _al_u852_o;
  wire _al_u853_o;
  wire _al_u854_o;
  wire _al_u855_o;
  wire _al_u856_o;
  wire _al_u857_o;
  wire _al_u859_o;
  wire _al_u860_o;
  wire _al_u861_o;
  wire _al_u862_o;
  wire _al_u863_o;
  wire _al_u864_o;
  wire _al_u865_o;
  wire _al_u866_o;
  wire _al_u867_o;
  wire _al_u868_o;
  wire _al_u869_o;
  wire _al_u870_o;
  wire _al_u871_o;
  wire _al_u872_o;
  wire _al_u873_o;
  wire _al_u874_o;
  wire _al_u875_o;
  wire _al_u876_o;
  wire _al_u877_o;
  wire _al_u878_o;
  wire _al_u880_o;
  wire _al_u881_o;
  wire _al_u882_o;
  wire _al_u883_o;
  wire _al_u884_o;
  wire _al_u885_o;
  wire _al_u886_o;
  wire _al_u887_o;
  wire _al_u888_o;
  wire _al_u889_o;
  wire _al_u890_o;
  wire _al_u891_o;
  wire _al_u892_o;
  wire _al_u893_o;
  wire _al_u894_o;
  wire _al_u895_o;
  wire _al_u896_o;
  wire _al_u897_o;
  wire _al_u898_o;
  wire _al_u899_o;
  wire _al_u901_o;
  wire _al_u902_o;
  wire _al_u903_o;
  wire _al_u904_o;
  wire _al_u905_o;
  wire _al_u906_o;
  wire _al_u907_o;
  wire _al_u908_o;
  wire _al_u909_o;
  wire _al_u910_o;
  wire _al_u911_o;
  wire _al_u912_o;
  wire _al_u913_o;
  wire _al_u914_o;
  wire _al_u915_o;
  wire _al_u916_o;
  wire _al_u917_o;
  wire _al_u918_o;
  wire _al_u919_o;
  wire _al_u920_o;
  wire _al_u922_o;
  wire _al_u923_o;
  wire _al_u924_o;
  wire _al_u925_o;
  wire _al_u926_o;
  wire _al_u927_o;
  wire _al_u928_o;
  wire _al_u929_o;
  wire _al_u930_o;
  wire _al_u931_o;
  wire _al_u932_o;
  wire _al_u933_o;
  wire _al_u934_o;
  wire _al_u935_o;
  wire _al_u936_o;
  wire _al_u937_o;
  wire _al_u938_o;
  wire _al_u939_o;
  wire _al_u940_o;
  wire _al_u941_o;
  wire _al_u943_o;
  wire _al_u944_o;
  wire _al_u945_o;
  wire _al_u946_o;
  wire _al_u947_o;
  wire _al_u948_o;
  wire _al_u949_o;
  wire _al_u950_o;
  wire _al_u951_o;
  wire _al_u952_o;
  wire _al_u953_o;
  wire _al_u954_o;
  wire _al_u955_o;
  wire _al_u956_o;
  wire _al_u957_o;
  wire _al_u958_o;
  wire _al_u959_o;
  wire _al_u960_o;
  wire _al_u961_o;
  wire _al_u962_o;
  wire _al_u964_o;
  wire _al_u965_o;
  wire _al_u966_o;
  wire _al_u967_o;
  wire _al_u968_o;
  wire _al_u969_o;
  wire _al_u970_o;
  wire _al_u971_o;
  wire _al_u972_o;
  wire _al_u973_o;
  wire _al_u974_o;
  wire _al_u975_o;
  wire _al_u976_o;
  wire _al_u977_o;
  wire _al_u978_o;
  wire _al_u979_o;
  wire _al_u980_o;
  wire _al_u981_o;
  wire _al_u982_o;
  wire _al_u983_o;
  wire _al_u985_o;
  wire _al_u986_o;
  wire _al_u987_o;
  wire _al_u988_o;
  wire _al_u989_o;
  wire _al_u990_o;
  wire _al_u991_o;
  wire _al_u992_o;
  wire _al_u993_o;
  wire _al_u994_o;
  wire _al_u995_o;
  wire _al_u996_o;
  wire _al_u997_o;
  wire _al_u998_o;
  wire _al_u999_o;
  wire clock_pad;  // __top.v(4)
  wire lt0_c1;
  wire lt0_c11;
  wire lt0_c13;
  wire lt0_c15;
  wire lt0_c17;
  wire lt0_c19;
  wire lt0_c21;
  wire lt0_c23;
  wire lt0_c25;
  wire lt0_c27;
  wire lt0_c29;
  wire lt0_c3;
  wire lt0_c31;
  wire lt0_c5;
  wire lt0_c7;
  wire lt0_c9;
  wire \m/dram_c0_mode ;
  wire \m/dram_c0_wclk ;
  wire \m/dram_c0_we ;
  wire \m/dram_c1_mode ;
  wire \m/dram_c1_wclk ;
  wire \m/dram_c1_we ;
  wire \m/dram_c2_mode ;
  wire \m/dram_c2_wclk ;
  wire \m/dram_c2_we ;
  wire \m/dram_c3_mode ;
  wire \m/dram_c3_wclk ;
  wire \m/dram_c3_we ;
  wire \m/dram_c4_mode ;
  wire \m/dram_c4_wclk ;
  wire \m/dram_c4_we ;
  wire \m/dram_c5_mode ;
  wire \m/dram_c5_wclk ;
  wire \m/dram_c5_we ;
  wire \m/dram_c6_mode ;
  wire \m/dram_c6_wclk ;
  wire \m/dram_c6_we ;
  wire \m/dram_c7_mode ;
  wire \m/dram_c7_wclk ;
  wire \m/dram_c7_we ;
  wire memwrite_cs;  // __top.v(14)
  wire n0;
  wire n7;
  wire rst_pad;  // __top.v(3)
  wire \t/a/WB_regwritecs ;  // cpu.v(69)
  wire \t/a/alu/add0/c11 ;
  wire \t/a/alu/add0/c15 ;
  wire \t/a/alu/add0/c19 ;
  wire \t/a/alu/add0/c23 ;
  wire \t/a/alu/add0/c27 ;
  wire \t/a/alu/add0/c3 ;
  wire \t/a/alu/add0/c31 ;
  wire \t/a/alu/add0/c7 ;
  wire \t/a/alu/lt0_c1 ;
  wire \t/a/alu/lt0_c11 ;
  wire \t/a/alu/lt0_c13 ;
  wire \t/a/alu/lt0_c15 ;
  wire \t/a/alu/lt0_c17 ;
  wire \t/a/alu/lt0_c19 ;
  wire \t/a/alu/lt0_c21 ;
  wire \t/a/alu/lt0_c23 ;
  wire \t/a/alu/lt0_c25 ;
  wire \t/a/alu/lt0_c27 ;
  wire \t/a/alu/lt0_c29 ;
  wire \t/a/alu/lt0_c3 ;
  wire \t/a/alu/lt0_c31 ;
  wire \t/a/alu/lt0_c5 ;
  wire \t/a/alu/lt0_c7 ;
  wire \t/a/alu/lt0_c9 ;
  wire \t/a/alu/n104_lutinv ;
  wire \t/a/alu/n105_lutinv ;
  wire \t/a/alu/n106_lutinv ;
  wire \t/a/alu/n132_lutinv ;
  wire \t/a/alu/n133_lutinv ;
  wire \t/a/alu/n134_lutinv ;
  wire \t/a/alu/n135_lutinv ;
  wire \t/a/alu/n136_lutinv ;
  wire \t/a/alu/n137_lutinv ;
  wire \t/a/alu/n138_lutinv ;
  wire \t/a/alu/n142_lutinv ;
  wire \t/a/alu/n143_lutinv ;
  wire \t/a/alu/n144_lutinv ;
  wire \t/a/alu/n145_lutinv ;
  wire \t/a/alu/n146_lutinv ;
  wire \t/a/alu/n147_lutinv ;
  wire \t/a/alu/n148_lutinv ;
  wire \t/a/alu/n149_lutinv ;
  wire \t/a/alu/n150_lutinv ;
  wire \t/a/alu/n151_lutinv ;
  wire \t/a/alu/n152_lutinv ;
  wire \t/a/alu/n153_lutinv ;
  wire \t/a/alu/n154_lutinv ;
  wire \t/a/alu/n155_lutinv ;
  wire \t/a/alu/n156_lutinv ;
  wire \t/a/alu/n157_lutinv ;
  wire \t/a/alu/n158_lutinv ;
  wire \t/a/alu/n159_lutinv ;
  wire \t/a/alu/n160_lutinv ;
  wire \t/a/alu/n161_lutinv ;
  wire \t/a/alu/n162_lutinv ;
  wire \t/a/alu/n163_lutinv ;
  wire \t/a/alu/n164_lutinv ;
  wire \t/a/alu/n165_lutinv ;
  wire \t/a/alu/n166_lutinv ;
  wire \t/a/alu/n167_lutinv ;
  wire \t/a/alu/n168_lutinv ;
  wire \t/a/alu/n169_lutinv ;
  wire \t/a/alu/n170_lutinv ;
  wire \t/a/alu/n173_lutinv ;
  wire \t/a/alu/n17_lutinv ;
  wire \t/a/alu/n18_lutinv ;
  wire \t/a/alu/n19_lutinv ;
  wire \t/a/alu/n202_lutinv ;
  wire \t/a/alu/n204_lutinv ;
  wire \t/a/alu/n20_lutinv ;
  wire \t/a/alu/n21_lutinv ;
  wire \t/a/alu/n22_lutinv ;
  wire \t/a/alu/n232_lutinv ;
  wire \t/a/alu/n233_lutinv ;
  wire \t/a/alu/n234_lutinv ;
  wire \t/a/alu/n23_lutinv ;
  wire \t/a/alu/n24_lutinv ;
  wire \t/a/alu/n25_lutinv ;
  wire \t/a/alu/n260_lutinv ;
  wire \t/a/alu/n261_lutinv ;
  wire \t/a/alu/n262_lutinv ;
  wire \t/a/alu/n263_lutinv ;
  wire \t/a/alu/n264_lutinv ;
  wire \t/a/alu/n265_lutinv ;
  wire \t/a/alu/n266_lutinv ;
  wire \t/a/alu/n26_lutinv ;
  wire \t/a/alu/n27_lutinv ;
  wire \t/a/alu/n28_lutinv ;
  wire \t/a/alu/n29_lutinv ;
  wire \t/a/alu/n30_lutinv ;
  wire \t/a/alu/n31_lutinv ;
  wire \t/a/alu/n32_lutinv ;
  wire \t/a/alu/n33_lutinv ;
  wire \t/a/alu/n34_lutinv ;
  wire \t/a/alu/n35_lutinv ;
  wire \t/a/alu/n36_lutinv ;
  wire \t/a/alu/n37_lutinv ;
  wire \t/a/alu/n38_lutinv ;
  wire \t/a/alu/n39_lutinv ;
  wire \t/a/alu/n40_lutinv ;
  wire \t/a/alu/n41_lutinv ;
  wire \t/a/alu/n42_lutinv ;
  wire \t/a/alu/n43_lutinv ;
  wire \t/a/alu/n44_lutinv ;
  wire \t/a/alu/n45_lutinv ;
  wire \t/a/alu/n56_lutinv ;
  wire \t/a/alu/n57_lutinv ;
  wire \t/a/alu/n8 ;
  wire \t/a/alu/sub0/c11 ;
  wire \t/a/alu/sub0/c15 ;
  wire \t/a/alu/sub0/c19 ;
  wire \t/a/alu/sub0/c23 ;
  wire \t/a/alu/sub0/c27 ;
  wire \t/a/alu/sub0/c3 ;
  wire \t/a/alu/sub0/c31 ;
  wire \t/a/alu/sub0/c7 ;
  wire \t/a/aluin/n10_lutinv ;
  wire \t/a/aluin/n11_lutinv ;
  wire \t/a/aluin/n12_lutinv ;
  wire \t/a/aluin/n35_lutinv ;
  wire \t/a/aluin/n5_lutinv ;
  wire \t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/condition/add0/c11 ;
  wire \t/a/condition/add0/c15 ;
  wire \t/a/condition/add0/c19 ;
  wire \t/a/condition/add0/c23 ;
  wire \t/a/condition/add0/c27 ;
  wire \t/a/condition/add0/c3 ;
  wire \t/a/condition/add0/c31 ;
  wire \t/a/condition/add0/c7 ;
  wire \t/a/condition/lt0_c1 ;
  wire \t/a/condition/lt0_c11 ;
  wire \t/a/condition/lt0_c13 ;
  wire \t/a/condition/lt0_c15 ;
  wire \t/a/condition/lt0_c17 ;
  wire \t/a/condition/lt0_c19 ;
  wire \t/a/condition/lt0_c21 ;
  wire \t/a/condition/lt0_c23 ;
  wire \t/a/condition/lt0_c25 ;
  wire \t/a/condition/lt0_c27 ;
  wire \t/a/condition/lt0_c29 ;
  wire \t/a/condition/lt0_c3 ;
  wire \t/a/condition/lt0_c31 ;
  wire \t/a/condition/lt0_c5 ;
  wire \t/a/condition/lt0_c7 ;
  wire \t/a/condition/lt0_c9 ;
  wire \t/a/condition/lt1_c1 ;
  wire \t/a/condition/lt1_c11 ;
  wire \t/a/condition/lt1_c13 ;
  wire \t/a/condition/lt1_c15 ;
  wire \t/a/condition/lt1_c17 ;
  wire \t/a/condition/lt1_c19 ;
  wire \t/a/condition/lt1_c21 ;
  wire \t/a/condition/lt1_c23 ;
  wire \t/a/condition/lt1_c25 ;
  wire \t/a/condition/lt1_c27 ;
  wire \t/a/condition/lt1_c29 ;
  wire \t/a/condition/lt1_c3 ;
  wire \t/a/condition/lt1_c31 ;
  wire \t/a/condition/lt1_c5 ;
  wire \t/a/condition/lt1_c7 ;
  wire \t/a/condition/lt1_c9 ;
  wire \t/a/condition/n0_lutinv ;
  wire \t/a/condition/n10 ;
  wire \t/a/condition/n1_lutinv ;
  wire \t/a/condition/n9 ;
  wire \t/a/ex_mem/n0 ;
  wire \t/a/if_id/n9 ;
  wire \t/a/instr/add0/c11 ;
  wire \t/a/instr/add0/c15 ;
  wire \t/a/instr/add0/c19 ;
  wire \t/a/instr/add0/c23 ;
  wire \t/a/instr/add0/c27 ;
  wire \t/a/instr/add0/c3 ;
  wire \t/a/instr/add0/c31 ;
  wire \t/a/instr/add0/c7 ;
  wire \t/a/instr/add2/c11 ;
  wire \t/a/instr/add2/c15 ;
  wire \t/a/instr/add2/c19 ;
  wire \t/a/instr/add2/c23 ;
  wire \t/a/instr/add2/c27 ;
  wire \t/a/instr/add2/c3 ;
  wire \t/a/instr/add2/c7 ;
  wire \t/a/n0_lutinv ;
  wire \t/a/n19 ;
  wire \t/a/n2 ;
  wire \t/a/n24_lutinv ;
  wire \t/a/n29 ;
  wire \t/a/n4_lutinv ;
  wire \t/a/n9_lutinv ;
  wire \t/a/regfile/mux39_b0_sel_is_3_o ;
  wire \t/a/regfile/mux39_b1000_sel_is_3_o ;
  wire \t/a/regfile/mux39_b100_sel_is_3_o ;
  wire \t/a/regfile/mux39_b128_sel_is_3_o ;
  wire \t/a/regfile/mux39_b160_sel_is_3_o ;
  wire \t/a/regfile/mux39_b192_sel_is_3_o ;
  wire \t/a/regfile/mux39_b224_sel_is_3_o ;
  wire \t/a/regfile/mux39_b256_sel_is_3_o ;
  wire \t/a/regfile/mux39_b288_sel_is_3_o ;
  wire \t/a/regfile/mux39_b320_sel_is_3_o ;
  wire \t/a/regfile/mux39_b32_sel_is_3_o ;
  wire \t/a/regfile/mux39_b352_sel_is_3_o ;
  wire \t/a/regfile/mux39_b384_sel_is_3_o ;
  wire \t/a/regfile/mux39_b416_sel_is_3_o ;
  wire \t/a/regfile/mux39_b448_sel_is_3_o ;
  wire \t/a/regfile/mux39_b480_sel_is_3_o ;
  wire \t/a/regfile/mux39_b512_sel_is_3_o ;
  wire \t/a/regfile/mux39_b544_sel_is_3_o ;
  wire \t/a/regfile/mux39_b576_sel_is_3_o ;
  wire \t/a/regfile/mux39_b608_sel_is_3_o ;
  wire \t/a/regfile/mux39_b640_sel_is_3_o ;
  wire \t/a/regfile/mux39_b64_sel_is_3_o ;
  wire \t/a/regfile/mux39_b672_sel_is_3_o ;
  wire \t/a/regfile/mux39_b704_sel_is_3_o ;
  wire \t/a/regfile/mux39_b736_sel_is_3_o ;
  wire \t/a/regfile/mux39_b768_sel_is_3_o ;
  wire \t/a/regfile/mux39_b800_sel_is_3_o ;
  wire \t/a/regfile/mux39_b832_sel_is_3_o ;
  wire \t/a/regfile/mux39_b864_sel_is_3_o ;
  wire \t/a/regfile/mux39_b896_sel_is_3_o ;
  wire \t/a/regfile/mux39_b928_sel_is_3_o ;
  wire \t/a/regfile/mux39_b960_sel_is_3_o ;
  wire \t/a/regfile/n1_lutinv ;
  wire \t/a/regfile/n3_lutinv ;
  wire \t/a/risk_jump/n11_lutinv ;
  wire \t/a/risk_jump/n19 ;
  wire \t/a/risk_jump/n24_lutinv ;
  wire \t/a/risk_jump/n35_lutinv ;
  wire \t/a/risk_jump/n42_lutinv ;
  wire \t/a/unconditional/eq1/or_xor_i0$5$_i1$5$_o_o_lutinv ;
  wire \t/busarbitration/mux5_b0_sel_is_3_o ;
  wire \t/busarbitration/mux6_b16_sel_is_3_o ;
  wire \t/busarbitration/n3 ;
  wire \t/instrnop ;  // top2.v(12)
  wire \t/instruction$2$_neg_lutinv ;
  wire \t/instruction$3$_neg_lutinv ;
  wire \t/instruction$4$_neg_lutinv ;
  wire \u1/c1 ;
  wire \u1/c11 ;
  wire \u1/c13 ;
  wire \u1/c15 ;
  wire \u1/c17 ;
  wire \u1/c19 ;
  wire \u1/c21 ;
  wire \u1/c23 ;
  wire \u1/c25 ;
  wire \u1/c27 ;
  wire \u1/c29 ;
  wire \u1/c3 ;
  wire \u1/c5 ;
  wire \u1/c7 ;
  wire \u1/c9 ;
  wire \u3/c11 ;
  wire \u3/c15 ;
  wire \u3/c19 ;
  wire \u3/c23 ;
  wire \u3/c27 ;
  wire \u3/c3 ;
  wire \u3/c7 ;

  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUT1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUT0(16'b0111000000110000),
    .INIT_LUT1(16'b1111000010110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1000 (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .d({\t/a/regfile/regfile$30$ [0],\t/a/regfile/regfile$30$ [0]}),
    .mi({open_n12,\t/a/regfile/regfile$31$ [0]}),
    .fx({open_n17,_al_u1000_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*B*A)"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(1*D*~C*B*A)"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1001|t/a/regfile/reg0_b928  (
    .a({_al_u1000_o,_al_u256_o}),
    .b({\t/a/ID_rs1 [0],\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$28$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$29$ [0],\t/a/WB_rd [3]}),
    .mi({open_n21,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1001_o,\t/a/regfile/mux39_b928_sel_is_3_o }),
    .q({open_n36,\t/a/regfile/regfile$29$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1002|_al_u1718  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs2 [2]}),
    .d({\t/a/regfile/regfile$26$ [0],\t/a/regfile/regfile$26$ [0]}),
    .e({\t/a/regfile/regfile$27$ [0],\t/a/regfile/regfile$27$ [0]}),
    .f({_al_u1002_o,_al_u1718_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1004|_al_u1003  (
    .a({_al_u999_o,_al_u1002_o}),
    .b({_al_u1001_o,\t/a/ID_rs1 [0]}),
    .c({_al_u1003_o,\t/a/ID_rs1 [1]}),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$24$ [0]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$25$ [0]}),
    .f({_al_u1004_o,_al_u1003_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*~(D*C))"),
    //.LUTF1("(~D*C*~B*A)"),
    //.LUTG0("(~1*B*A*~(D*C))"),
    //.LUTG1("(~D*C*~B*A)"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0000000000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1006|_al_u1038  (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_fun3 [0],\t/a/MEM_regdat2 [0]}),
    .c(\t/a/MEM_fun3 [1:0]),
    .d(\t/a/MEM_fun3 [2:1]),
    .e({open_n83,\t/a/MEM_fun3 [2]}),
    .f({\t/busarbitration/mux6_b16_sel_is_3_o ,o_data[0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1007|_al_u1022  (
    .c({\t/a/MEM_regdat2 [31],\t/a/MEM_regdat2 [16]}),
    .d({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .f({o_data[31],o_data[16]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1008|_al_u1021  (
    .c({\t/a/MEM_regdat2 [30],\t/a/MEM_regdat2 [17]}),
    .d({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .f({o_data[30],o_data[17]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1009|_al_u1020  (
    .c({\t/a/MEM_regdat2 [29],\t/a/MEM_regdat2 [18]}),
    .d({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .f({o_data[29],o_data[18]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1010|_al_u1019  (
    .c({\t/a/MEM_regdat2 [28],\t/a/MEM_regdat2 [19]}),
    .d({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .f({o_data[28],o_data[19]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1011|_al_u1018  (
    .c({\t/a/MEM_regdat2 [27],\t/a/MEM_regdat2 [20]}),
    .d({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .f({o_data[27],o_data[20]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1012|_al_u1017  (
    .c({\t/a/MEM_regdat2 [26],\t/a/MEM_regdat2 [21]}),
    .d({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .f({o_data[26],o_data[21]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1013|_al_u1016  (
    .c({\t/a/MEM_regdat2 [25],\t/a/MEM_regdat2 [22]}),
    .d({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .f({o_data[25],o_data[22]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1014|_al_u1015  (
    .c(\t/a/MEM_regdat2 [24:23]),
    .d({\t/busarbitration/mux6_b16_sel_is_3_o ,\t/busarbitration/mux6_b16_sel_is_3_o }),
    .f(o_data[24:23]));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*~(D*C))"),
    //.LUTF1("(~0*B*A*(D@C))"),
    //.LUTG0("(~1*B*A*~(D*C))"),
    //.LUTG1("(~1*B*A*(D@C))"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0000100010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1023|_al_u1035  (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [9],\t/a/MEM_regdat2 [3]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .e({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [2]}),
    .f({o_data[9],o_data[3]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*~(D*C))"),
    //.LUTF1("(~0*B*A*(D@C))"),
    //.LUTG0("(~1*B*A*~(D*C))"),
    //.LUTG1("(~1*B*A*(D@C))"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0000100010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1024|_al_u1034  (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [8],\t/a/MEM_regdat2 [4]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .e({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [2]}),
    .f({o_data[8],o_data[4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*~(D*C))"),
    //.LUTF1("(~0*B*A*(D@C))"),
    //.LUTG0("(~1*B*A*~(D*C))"),
    //.LUTG1("(~1*B*A*(D@C))"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0000100010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1025|_al_u1031  (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [15],\t/a/MEM_regdat2 [7]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .e({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [2]}),
    .f({o_data[15],o_data[7]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*(D@C))"),
    //.LUTF1("(~0*B*A*(D@C))"),
    //.LUTG0("(~1*B*A*(D@C))"),
    //.LUTG1("(~1*B*A*(D@C))"),
    .INIT_LUTF0(16'b0000100010000000),
    .INIT_LUTF1(16'b0000100010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1026|_al_u1030  (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [14],\t/a/MEM_regdat2 [10]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .e({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [2]}),
    .f({o_data[14],o_data[10]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*(D@C))"),
    //.LUT1("(~1*B*A*(D@C))"),
    .INIT_LUT0(16'b0000100010000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1028 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [12],\t/a/MEM_regdat2 [12]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .mi({open_n412,\t/a/MEM_fun3 [2]}),
    .fx({open_n417,o_data[12]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*(D@C))"),
    //.LUT1("(~1*B*A*(D@C))"),
    .INIT_LUT0(16'b0000100010000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1029 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [11],\t/a/MEM_regdat2 [11]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .mi({open_n432,\t/a/MEM_fun3 [2]}),
    .fx({open_n437,o_data[11]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*~(D*C))"),
    //.LUT1("(~1*B*A*~(D*C))"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1032 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [6],\t/a/MEM_regdat2 [6]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .mi({open_n452,\t/a/MEM_fun3 [2]}),
    .fx({open_n457,o_data[6]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*~(D*C))"),
    //.LUT1("(~1*B*A*~(D*C))"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1033 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [5],\t/a/MEM_regdat2 [5]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .mi({open_n472,\t/a/MEM_fun3 [2]}),
    .fx({open_n477,o_data[5]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*~(D*C))"),
    //.LUT1("(~1*B*A*~(D*C))"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1036 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [2],\t/a/MEM_regdat2 [2]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .mi({open_n492,\t/a/MEM_fun3 [2]}),
    .fx({open_n497,o_data[2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*B*A*~(D*C))"),
    //.LUT1("(~1*B*A*~(D*C))"),
    .INIT_LUT0(16'b0000100010001000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1037 (
    .a({memwrite_cs,memwrite_cs}),
    .b({\t/a/MEM_regdat2 [1],\t/a/MEM_regdat2 [1]}),
    .c({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [0]}),
    .d({\t/a/MEM_fun3 [1],\t/a/MEM_fun3 [1]}),
    .mi({open_n512,\t/a/MEM_fun3 [2]}),
    .fx({open_n517,o_data[1]}));
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1039|t/a/if_id/reg5_b5  (
    .b({open_n522,\t/a/MEM_aludat [5]}),
    .c({memwrite_cs,\t/memstraddress [5]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[5],\t/busarbitration/n3 }),
    .mi({open_n533,\t/memstraddress [5]}),
    .sr(rst_pad),
    .f({n3[3],addr[5]}),
    .q({open_n537,\t/a/ID_memstraddr [5]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1040|_al_u297  (
    .b({open_n540,\t/a/MEM_aludat [4]}),
    .c({memwrite_cs,\t/memstraddress [4]}),
    .d({addr[4],\t/busarbitration/n3 }),
    .f({n3[2],addr[4]}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u1041|_al_u300  (
    .b({open_n563,\t/a/MEM_aludat [3]}),
    .c({memwrite_cs,\t/memstraddress [3]}),
    .d({addr[3],\t/busarbitration/n3 }),
    .f({n3[1],addr[3]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1042|_al_u311  (
    .b({open_n586,\t/a/MEM_aludat [2]}),
    .c({memwrite_cs,\t/memstraddress [2]}),
    .d({addr[2],\t/busarbitration/n3 }),
    .f({n3[0],addr[2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0@C)*~(D*~B))"),
    //.LUT1("(~A*~(1@C)*~(D*~B))"),
    .INIT_LUT0(16'b0000010000000101),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1044 (
    .a({_al_u1043_o,_al_u1043_o}),
    .b({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .c({\t/a/ID_rs2 [4],\t/a/ID_rs2 [4]}),
    .d({\t/a/WB_rd [2],\t/a/WB_rd [2]}),
    .mi({open_n623,\t/a/WB_rd [4]}),
    .fx({open_n628,_al_u1044_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~0*C)*~(D*~B))"),
    //.LUT1("(A*~(~1*C)*~(D*~B))"),
    .INIT_LUT0(16'b0000100000001010),
    .INIT_LUT1(16'b1000100010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1045 (
    .a({_al_u1044_o,_al_u1044_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .d({\t/a/WB_rd [0],\t/a/WB_rd [0]}),
    .mi({open_n643,\t/a/WB_rd [2]}),
    .fx({open_n648,_al_u1045_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1048|_al_u1047  (
    .a({open_n651,_al_u1046_o}),
    .b({open_n652,\t/a/ID_rs2 [1]}),
    .c({_al_u1047_o,\t/a/ID_rs2 [3]}),
    .d({_al_u1045_o,\t/a/WB_rd [1]}),
    .e({open_n655,\t/a/WB_rd [3]}),
    .f({\t/a/regfile/n3_lutinv ,_al_u1047_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*~B*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(1*D*~C*~B*A)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1049|_al_u2604  (
    .a({open_n676,\t/a/regfile/n3_lutinv }),
    .b({open_n677,\t/a/risk_jump/n42_lutinv }),
    .c({\t/a/WB_regwritecs ,\t/a/risk_jump/n35_lutinv }),
    .d({\t/a/regfile/n3_lutinv ,\t/a/n19 }),
    .e({open_n680,\t/a/condition/n1_lutinv }),
    .f({_al_u1049_o,_al_u2604_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1050|_al_u1505  (
    .a({\t/a/ID_rs2 [0],_al_u1501_o}),
    .b({\t/a/ID_rs2 [1],_al_u1502_o}),
    .c({\t/a/regfile/regfile$4$ [9],_al_u1503_o}),
    .d({\t/a/regfile/regfile$5$ [9],_al_u1504_o}),
    .e({open_n703,\t/a/ID_rs2 [2]}),
    .f({_al_u1050_o,_al_u1505_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1053|t/a/regfile/reg0_b73  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [9],\t/a/regfile/regfile$3$ [9]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [9],\t/a/regfile/regfile$2$ [9]}),
    .mi({open_n734,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u1053_o,_al_u347_o}),
    .q({open_n738,\t/a/regfile/regfile$2$ [9]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1054 (
    .a({_al_u1050_o,_al_u1050_o}),
    .b({_al_u1051_o,_al_u1051_o}),
    .c({_al_u1052_o,_al_u1052_o}),
    .d({_al_u1053_o,_al_u1053_o}),
    .mi({open_n751,\t/a/ID_rs2 [2]}),
    .fx({open_n756,_al_u1054_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1059|t/a/regfile/reg0_b425  (
    .a({_al_u1054_o,_al_u1055_o}),
    .b({_al_u1056_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1058_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [9]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [9]}),
    .mi({open_n760,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u1059_o,_al_u1056_o}),
    .q({open_n775,\t/a/regfile/regfile$13$ [9]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1064 (
    .a({_al_u1060_o,_al_u1060_o}),
    .b({_al_u1061_o,_al_u1061_o}),
    .c({_al_u1062_o,_al_u1062_o}),
    .d({_al_u1063_o,_al_u1063_o}),
    .mi({open_n788,\t/a/ID_rs2 [2]}),
    .fx({open_n793,_al_u1064_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1069|t/a/regfile/reg0_b937  (
    .a({_al_u1064_o,_al_u1065_o}),
    .b({_al_u1066_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1068_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [9]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [9]}),
    .mi({open_n797,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u1069_o,_al_u1066_o}),
    .q({open_n812,\t/a/regfile/regfile$29$ [9]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1072|t/a/regfile/reg0_b968  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [8],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [8],\t/a/regfile/regfile$31$ [8]}),
    .e({open_n813,\t/a/regfile/regfile$30$ [8]}),
    .mi({open_n815,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u1072_o,_al_u370_o}),
    .q({open_n830,\t/a/regfile/regfile$30$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1075|_al_u1285  (
    .a({_al_u1071_o,_al_u1281_o}),
    .b({_al_u1072_o,_al_u1282_o}),
    .c({_al_u1073_o,_al_u1283_o}),
    .d({_al_u1074_o,_al_u1284_o}),
    .e({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .f({_al_u1075_o,_al_u1285_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1080|t/a/regfile/reg0_b680  (
    .a({_al_u1075_o,_al_u1076_o}),
    .b({_al_u1077_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1079_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$20$ [8]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [8]}),
    .mi({open_n854,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u1080_o,_al_u1077_o}),
    .q({open_n869,\t/a/regfile/regfile$21$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1081|_al_u1327  (
    .a({\t/a/ID_rs2 [0],_al_u1323_o}),
    .b({\t/a/ID_rs2 [1],_al_u1324_o}),
    .c({\t/a/regfile/regfile$4$ [8],_al_u1325_o}),
    .d({\t/a/regfile/regfile$5$ [8],_al_u1326_o}),
    .e({open_n872,\t/a/ID_rs2 [2]}),
    .f({_al_u1081_o,_al_u1327_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1082|_al_u1369  (
    .a({\t/a/ID_rs2 [0],_al_u1365_o}),
    .b({\t/a/ID_rs2 [1],_al_u1366_o}),
    .c({\t/a/regfile/regfile$6$ [8],_al_u1367_o}),
    .d({\t/a/regfile/regfile$7$ [8],_al_u1368_o}),
    .e({open_n895,\t/a/ID_rs2 [2]}),
    .f({_al_u1082_o,_al_u1369_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1084|t/a/regfile/reg0_b72  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [8],\t/a/regfile/regfile$3$ [8]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [8],\t/a/regfile/regfile$2$ [8]}),
    .mi({open_n926,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u1084_o,_al_u358_o}),
    .q({open_n930,\t/a/regfile/regfile$2$ [8]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1090|t/a/regfile/reg0_b424  (
    .a({_al_u1085_o,_al_u1086_o}),
    .b({_al_u1087_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1089_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [8]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [8]}),
    .mi({open_n932,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u1090_o,_al_u1087_o}),
    .q({open_n947,\t/a/regfile/regfile$13$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1092|_al_u1096  (
    .a({\t/a/ID_rs2 [0],_al_u1092_o}),
    .b({\t/a/ID_rs2 [1],_al_u1093_o}),
    .c({\t/a/regfile/regfile$4$ [7],_al_u1094_o}),
    .d({\t/a/regfile/regfile$5$ [7],_al_u1095_o}),
    .e({open_n950,\t/a/ID_rs2 [2]}),
    .f({_al_u1092_o,_al_u1096_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1095|t/a/regfile/reg0_b71  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [7],\t/a/regfile/regfile$3$ [7]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [7],\t/a/regfile/regfile$2$ [7]}),
    .mi({open_n981,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({_al_u1095_o,_al_u389_o}),
    .q({open_n985,\t/a/regfile/regfile$2$ [7]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1101|t/a/regfile/reg0_b423  (
    .a({_al_u1096_o,_al_u1097_o}),
    .b({_al_u1098_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1100_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [7]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [7]}),
    .mi({open_n987,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({_al_u1101_o,_al_u1098_o}),
    .q({open_n1002,\t/a/regfile/regfile$13$ [7]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1106|_al_u1421  (
    .a({_al_u1102_o,_al_u1417_o}),
    .b({_al_u1103_o,_al_u1418_o}),
    .c({_al_u1104_o,_al_u1419_o}),
    .d({_al_u1105_o,_al_u1420_o}),
    .e({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .f({_al_u1106_o,_al_u1421_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1111|t/a/regfile/reg0_b935  (
    .a({_al_u1106_o,_al_u1107_o}),
    .b({_al_u1108_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1110_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [7]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [7]}),
    .mi({open_n1026,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({_al_u1111_o,_al_u1108_o}),
    .q({open_n1041,\t/a/regfile/regfile$29$ [7]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1113|t/a/regfile/reg0_b134  (
    .a({\t/a/ID_rs2 [0],_al_u2606_o}),
    .b({\t/a/ID_rs2 [1],_al_u2610_o}),
    .c({\t/a/regfile/regfile$4$ [6],\t/a/MEM_aludat [6]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [6],\t/a/reg_writedat [6]}),
    .mi({open_n1052,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u1113_o,_al_u2730_o}),
    .q({open_n1056,\t/a/regfile/regfile$4$ [6]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1116|t/a/regfile/reg0_b70  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [6],\t/a/regfile/regfile$3$ [6]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [6],\t/a/regfile/regfile$2$ [6]}),
    .mi({open_n1067,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u1116_o,_al_u400_o}),
    .q({open_n1071,\t/a/regfile/regfile$2$ [6]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1117 (
    .a({_al_u1113_o,_al_u1113_o}),
    .b({_al_u1114_o,_al_u1114_o}),
    .c({_al_u1115_o,_al_u1115_o}),
    .d({_al_u1116_o,_al_u1116_o}),
    .mi({open_n1084,\t/a/ID_rs2 [2]}),
    .fx({open_n1089,_al_u1117_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1122|t/a/regfile/reg0_b422  (
    .a({_al_u1117_o,_al_u1118_o}),
    .b({_al_u1119_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1121_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [6]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [6]}),
    .mi({open_n1093,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u1122_o,_al_u1119_o}),
    .q({open_n1108,\t/a/regfile/regfile$13$ [6]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1127 (
    .a({_al_u1123_o,_al_u1123_o}),
    .b({_al_u1124_o,_al_u1124_o}),
    .c({_al_u1125_o,_al_u1125_o}),
    .d({_al_u1126_o,_al_u1126_o}),
    .mi({open_n1121,\t/a/ID_rs2 [2]}),
    .fx({open_n1126,_al_u1127_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1132|t/a/regfile/reg0_b934  (
    .a({_al_u1127_o,_al_u1128_o}),
    .b({_al_u1129_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1131_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [6]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [6]}),
    .mi({open_n1130,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u1132_o,_al_u1129_o}),
    .q({open_n1145,\t/a/regfile/regfile$29$ [6]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1134|t/a/regfile/reg0_b133  (
    .a({\t/a/ID_rs2 [0],_al_u2606_o}),
    .b({\t/a/ID_rs2 [1],_al_u2610_o}),
    .c({\t/a/regfile/regfile$4$ [5],\t/a/MEM_aludat [5]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [5],\t/a/reg_writedat [5]}),
    .mi({open_n1156,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u1134_o,_al_u2737_o}),
    .q({open_n1160,\t/a/regfile/regfile$4$ [5]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1135|_al_u1138  (
    .a({\t/a/ID_rs2 [0],_al_u1134_o}),
    .b({\t/a/ID_rs2 [1],_al_u1135_o}),
    .c({\t/a/regfile/regfile$6$ [5],_al_u1136_o}),
    .d({\t/a/regfile/regfile$7$ [5],_al_u1137_o}),
    .e({open_n1163,\t/a/ID_rs2 [2]}),
    .f({_al_u1135_o,_al_u1138_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1137|t/a/regfile/reg0_b69  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [5],\t/a/regfile/regfile$3$ [5]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [5],\t/a/regfile/regfile$2$ [5]}),
    .mi({open_n1194,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u1137_o,_al_u421_o}),
    .q({open_n1198,\t/a/regfile/regfile$2$ [5]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1143|t/a/regfile/reg0_b421  (
    .a({_al_u1138_o,_al_u1139_o}),
    .b({_al_u1140_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1142_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [5]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [5]}),
    .mi({open_n1200,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u1143_o,_al_u1140_o}),
    .q({open_n1215,\t/a/regfile/regfile$13$ [5]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1148|_al_u1358  (
    .a({_al_u1144_o,_al_u1354_o}),
    .b({_al_u1145_o,_al_u1355_o}),
    .c({_al_u1146_o,_al_u1356_o}),
    .d({_al_u1147_o,_al_u1357_o}),
    .e({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .f({_al_u1148_o,_al_u1358_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1153|t/a/regfile/reg0_b933  (
    .a({_al_u1148_o,_al_u1149_o}),
    .b({_al_u1150_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1152_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [5]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [5]}),
    .mi({open_n1239,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u1153_o,_al_u1150_o}),
    .q({open_n1254,\t/a/regfile/regfile$29$ [5]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1155|t/a/regfile/reg0_b164  (
    .a({\t/a/ID_rs2 [0],_al_u2606_o}),
    .b({\t/a/ID_rs2 [1],_al_u2610_o}),
    .c({\t/a/regfile/regfile$4$ [4],\t/a/MEM_aludat [4]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [4],\t/a/reg_writedat [4]}),
    .mi({open_n1265,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u1155_o,_al_u2742_o}),
    .q({open_n1269,\t/a/regfile/regfile$5$ [4]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~A*~(~0*B)))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(C*~(D*~A*~(~1*B)))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0101111100001111),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1156|t/a/regfile/reg0_b196  (
    .a({\t/a/ID_rs2 [0],_al_u1999_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$6$ [4],_al_u2000_o}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [4],\t/a/aluin/n10_lutinv }),
    .e({open_n1270,\t/a/reg_writedat [4]}),
    .mi({open_n1272,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u1156_o,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .q({open_n1287,\t/a/regfile/regfile$6$ [4]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*C*B*A)"),
    //.LUTF1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(~1*~D*C*B*A)"),
    //.LUTG1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1158|t/a/regfile/reg0_b100  (
    .a({\t/a/ID_rs2 [0],_al_u254_o}),
    .b({\t/a/ID_rs2 [1],\t/a/WB_rd [0]}),
    .c({\t/a/regfile/regfile$3$ [4],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [4],\t/a/WB_rd [2]}),
    .e({open_n1288,\t/a/WB_rd [3]}),
    .mi({open_n1290,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u1158_o,\t/a/regfile/mux39_b100_sel_is_3_o }),
    .q({open_n1305,\t/a/regfile/regfile$3$ [4]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1164|t/a/regfile/reg0_b420  (
    .a({_al_u1159_o,_al_u1160_o}),
    .b({_al_u1161_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1163_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [4]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [4]}),
    .mi({open_n1307,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u1164_o,_al_u1161_o}),
    .q({open_n1322,\t/a/regfile/regfile$13$ [4]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1169|_al_u1316  (
    .a({_al_u1165_o,_al_u1312_o}),
    .b({_al_u1166_o,_al_u1313_o}),
    .c({_al_u1167_o,_al_u1314_o}),
    .d({_al_u1168_o,_al_u1315_o}),
    .e({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .f({_al_u1169_o,_al_u1316_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1174|t/a/regfile/reg0_b932  (
    .a({_al_u1169_o,_al_u1170_o}),
    .b({_al_u1171_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1173_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [4]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [4]}),
    .mi({open_n1346,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u1174_o,_al_u1171_o}),
    .q({open_n1361,\t/a/regfile/regfile$29$ [4]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1180|_al_u1222  (
    .a({_al_u1176_o,_al_u1218_o}),
    .b({_al_u1177_o,_al_u1219_o}),
    .c({_al_u1178_o,_al_u1220_o}),
    .d({_al_u1179_o,_al_u1221_o}),
    .e({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .f({_al_u1180_o,_al_u1222_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1185|t/a/regfile/reg0_b675  (
    .a({_al_u1180_o,_al_u1181_o}),
    .b({_al_u1182_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1184_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$20$ [3]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [3]}),
    .mi({open_n1385,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u1185_o,_al_u1182_o}),
    .q({open_n1400,\t/a/regfile/regfile$21$ [3]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1186|t/a/regfile/reg0_b131  (
    .a({\t/a/ID_rs2 [0],_al_u2614_o}),
    .b({\t/a/ID_rs2 [1],_al_u2616_o}),
    .c({\t/a/regfile/regfile$4$ [3],\t/a/MEM_aludat [3]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [3],\t/a/reg_writedat [3]}),
    .mi({open_n1411,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u1186_o,_al_u2752_o}),
    .q({open_n1415,\t/a/regfile/regfile$4$ [3]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~A*~(~0*B)))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(C*~(D*~A*~(~1*B)))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0101111100001111),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1187|t/a/regfile/reg0_b195  (
    .a({\t/a/ID_rs2 [0],_al_u2009_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$6$ [3],_al_u2010_o}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [3],\t/a/aluin/n10_lutinv }),
    .e({open_n1416,\t/a/reg_writedat [3]}),
    .mi({open_n1418,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u1187_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .q({open_n1433,\t/a/regfile/regfile$6$ [3]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1190 (
    .a({_al_u1186_o,_al_u1186_o}),
    .b({_al_u1187_o,_al_u1187_o}),
    .c({_al_u1188_o,_al_u1188_o}),
    .d({_al_u1189_o,_al_u1189_o}),
    .mi({open_n1446,\t/a/ID_rs2 [2]}),
    .fx({open_n1451,_al_u1190_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1195|t/a/regfile/reg0_b419  (
    .a({_al_u1190_o,_al_u1191_o}),
    .b({_al_u1192_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1194_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [3]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [3]}),
    .mi({open_n1455,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u1195_o,_al_u1192_o}),
    .q({open_n1470,\t/a/regfile/regfile$13$ [3]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1197|t/a/regfile/reg0_b191  (
    .a({\t/a/ID_rs2 [0],_al_u1823_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_A_select [1]}),
    .c({\t/a/regfile/regfile$4$ [31],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [31],\t/a/reg_writedat [31]}),
    .mi({open_n1474,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1197_o,\t/a/aluin/sel0_b31/B0 }),
    .q({open_n1489,\t/a/regfile/regfile$5$ [31]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1200|t/a/regfile/reg0_b95  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [31],\t/a/regfile/regfile$3$ [31]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [31],\t/a/regfile/regfile$2$ [31]}),
    .mi({open_n1500,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1200_o,_al_u494_o}),
    .q({open_n1504,\t/a/regfile/regfile$2$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1201 (
    .a({_al_u1197_o,_al_u1197_o}),
    .b({_al_u1198_o,_al_u1198_o}),
    .c({_al_u1199_o,_al_u1199_o}),
    .d({_al_u1200_o,_al_u1200_o}),
    .mi({open_n1517,\t/a/ID_rs2 [2]}),
    .fx({open_n1522,_al_u1201_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1206|t/a/regfile/reg0_b447  (
    .a({_al_u1201_o,_al_u1202_o}),
    .b({_al_u1203_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1205_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [31]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [31]}),
    .mi({open_n1526,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1206_o,_al_u1203_o}),
    .q({open_n1541,\t/a/regfile/regfile$13$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1211|_al_u1212  (
    .a({_al_u1207_o,\t/a/ID_rs2 [0]}),
    .b({_al_u1208_o,\t/a/ID_rs2 [1]}),
    .c({_al_u1209_o,\t/a/ID_rs2 [2]}),
    .d({_al_u1210_o,\t/a/regfile/regfile$31$ [31]}),
    .e({\t/a/ID_rs2 [2],\t/a/regfile/regfile$30$ [31]}),
    .f({_al_u1211_o,_al_u1212_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1216|t/a/regfile/reg0_b959  (
    .a({_al_u1211_o,_al_u1212_o}),
    .b({_al_u1213_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1215_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [31]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [31]}),
    .mi({open_n1565,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1216_o,_al_u1213_o}),
    .q({open_n1580,\t/a/regfile/regfile$29$ [31]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1219|t/a/regfile/reg0_b990  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [30],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [30],\t/a/regfile/regfile$31$ [30]}),
    .e({open_n1581,\t/a/regfile/regfile$30$ [30]}),
    .mi({open_n1583,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1219_o,_al_u517_o}),
    .q({open_n1598,\t/a/regfile/regfile$30$ [30]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1227|t/a/regfile/reg0_b702  (
    .a({_al_u1222_o,_al_u1223_o}),
    .b({_al_u1224_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1226_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$20$ [30]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [30]}),
    .mi({open_n1600,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1227_o,_al_u1224_o}),
    .q({open_n1615,\t/a/regfile/regfile$21$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1228|_al_u1232  (
    .a({\t/a/ID_rs2 [0],_al_u1228_o}),
    .b({\t/a/ID_rs2 [1],_al_u1229_o}),
    .c({\t/a/regfile/regfile$4$ [30],_al_u1230_o}),
    .d({\t/a/regfile/regfile$5$ [30],_al_u1231_o}),
    .e({open_n1618,\t/a/ID_rs2 [2]}),
    .f({_al_u1228_o,_al_u1232_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1231|t/a/regfile/reg0_b94  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [30],\t/a/regfile/regfile$3$ [30]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [30],\t/a/regfile/regfile$2$ [30]}),
    .mi({open_n1649,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1231_o,_al_u505_o}),
    .q({open_n1653,\t/a/regfile/regfile$2$ [30]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1237|t/a/regfile/reg0_b446  (
    .a({_al_u1232_o,_al_u1233_o}),
    .b({_al_u1234_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1236_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [30]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [30]}),
    .mi({open_n1655,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1237_o,_al_u1234_o}),
    .q({open_n1670,\t/a/regfile/regfile$13$ [30]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1239|t/a/regfile/reg0_b130  (
    .a({\t/a/ID_rs2 [0],_al_u2614_o}),
    .b({\t/a/ID_rs2 [1],_al_u2616_o}),
    .c({\t/a/regfile/regfile$4$ [2],\t/a/MEM_aludat [2]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [2],\t/a/reg_writedat [2]}),
    .mi({open_n1681,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u1239_o,_al_u2756_o}),
    .q({open_n1685,\t/a/regfile/regfile$4$ [2]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*(~A*~(0)*~(B)+~A*0*~(B)+~(~A)*0*B+~A*0*B)))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(C*~(D*(~A*~(1)*~(B)+~A*1*~(B)+~(~A)*1*B+~A*1*B)))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b1101111100001111),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1240|t/a/regfile/reg0_b194  (
    .a({\t/a/ID_rs2 [0],_al_u2092_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$6$ [2],_al_u2093_o}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [2],\t/a/aluin/n10_lutinv }),
    .e({open_n1686,\t/a/reg_writedat [2]}),
    .mi({open_n1688,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u1240_o,\t/a/EX_B [2]}),
    .q({open_n1703,\t/a/regfile/regfile$6$ [2]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1243 (
    .a({_al_u1239_o,_al_u1239_o}),
    .b({_al_u1240_o,_al_u1240_o}),
    .c({_al_u1241_o,_al_u1241_o}),
    .d({_al_u1242_o,_al_u1242_o}),
    .mi({open_n1716,\t/a/ID_rs2 [2]}),
    .fx({open_n1721,_al_u1243_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1248|t/a/regfile/reg0_b418  (
    .a({_al_u1243_o,_al_u1244_o}),
    .b({_al_u1245_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1247_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [2]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [2]}),
    .mi({open_n1725,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u1248_o,_al_u1245_o}),
    .q({open_n1740,\t/a/regfile/regfile$13$ [2]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1253|_al_u1274  (
    .a({_al_u1249_o,_al_u1270_o}),
    .b({_al_u1250_o,_al_u1271_o}),
    .c({_al_u1251_o,_al_u1272_o}),
    .d({_al_u1252_o,_al_u1273_o}),
    .e({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .f({_al_u1253_o,_al_u1274_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1258|t/a/regfile/reg0_b930  (
    .a({_al_u1253_o,_al_u1254_o}),
    .b({_al_u1255_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1257_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [2]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [2]}),
    .mi({open_n1764,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u1258_o,_al_u1255_o}),
    .q({open_n1779,\t/a/regfile/regfile$29$ [2]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1263|t/a/regfile/reg0_b93  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [29],\t/a/regfile/regfile$3$ [29]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [29],\t/a/regfile/regfile$2$ [29]}),
    .mi({open_n1790,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1263_o,_al_u557_o}),
    .q({open_n1794,\t/a/regfile/regfile$2$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1264 (
    .a({_al_u1260_o,_al_u1260_o}),
    .b({_al_u1261_o,_al_u1261_o}),
    .c({_al_u1262_o,_al_u1262_o}),
    .d({_al_u1263_o,_al_u1263_o}),
    .mi({open_n1807,\t/a/ID_rs2 [2]}),
    .fx({open_n1812,_al_u1264_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1269|t/a/regfile/reg0_b445  (
    .a({_al_u1264_o,_al_u1265_o}),
    .b({_al_u1266_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1268_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [29]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [29]}),
    .mi({open_n1816,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1269_o,_al_u1266_o}),
    .q({open_n1831,\t/a/regfile/regfile$13$ [29]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUT1("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .INIT_LUT0(16'b1011000000110000),
    .INIT_LUT1(16'b1111000001110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1275 (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .d({\t/a/regfile/regfile$31$ [29],\t/a/regfile/regfile$31$ [29]}),
    .mi({open_n1844,\t/a/regfile/regfile$30$ [29]}),
    .fx({open_n1849,_al_u1275_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1279|t/a/regfile/reg0_b957  (
    .a({_al_u1274_o,_al_u1275_o}),
    .b({_al_u1276_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1278_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [29]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [29]}),
    .mi({open_n1853,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1279_o,_al_u1276_o}),
    .q({open_n1868,\t/a/regfile/regfile$29$ [29]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1282|t/a/regfile/reg0_b988  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [28],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [28],\t/a/regfile/regfile$31$ [28]}),
    .e({open_n1869,\t/a/regfile/regfile$30$ [28]}),
    .mi({open_n1871,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1282_o,_al_u580_o}),
    .q({open_n1886,\t/a/regfile/regfile$30$ [28]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1290|t/a/regfile/reg0_b700  (
    .a({_al_u1285_o,_al_u1286_o}),
    .b({_al_u1287_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1289_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$20$ [28]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [28]}),
    .mi({open_n1888,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1290_o,_al_u1287_o}),
    .q({open_n1903,\t/a/regfile/regfile$21$ [28]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1291|t/a/regfile/reg0_b188  (
    .a({\t/a/ID_rs2 [0],_al_u1835_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_A_select [1]}),
    .c({\t/a/regfile/regfile$4$ [28],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [28],\t/a/reg_writedat [28]}),
    .mi({open_n1907,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1291_o,\t/a/aluin/sel0_b28/B0 }),
    .q({open_n1922,\t/a/regfile/regfile$5$ [28]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1294|t/a/regfile/reg0_b92  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [28],\t/a/regfile/regfile$3$ [28]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [28],\t/a/regfile/regfile$2$ [28]}),
    .mi({open_n1933,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1294_o,_al_u568_o}),
    .q({open_n1937,\t/a/regfile/regfile$2$ [28]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1295 (
    .a({_al_u1291_o,_al_u1291_o}),
    .b({_al_u1292_o,_al_u1292_o}),
    .c({_al_u1293_o,_al_u1293_o}),
    .d({_al_u1294_o,_al_u1294_o}),
    .mi({open_n1950,\t/a/ID_rs2 [2]}),
    .fx({open_n1955,_al_u1295_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1300|t/a/regfile/reg0_b444  (
    .a({_al_u1295_o,_al_u1296_o}),
    .b({_al_u1297_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1299_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [28]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [28]}),
    .mi({open_n1959,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1300_o,_al_u1297_o}),
    .q({open_n1974,\t/a/regfile/regfile$13$ [28]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1302|t/a/regfile/reg0_b187  (
    .a({\t/a/ID_rs2 [0],_al_u1838_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_A_select [1]}),
    .c({\t/a/regfile/regfile$4$ [27],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [27],\t/a/reg_writedat [27]}),
    .mi({open_n1978,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1302_o,\t/a/aluin/sel0_b27/B0 }),
    .q({open_n1993,\t/a/regfile/regfile$5$ [27]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1305|t/a/regfile/reg0_b91  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [27],\t/a/regfile/regfile$3$ [27]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [27],\t/a/regfile/regfile$2$ [27]}),
    .mi({open_n2004,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1305_o,_al_u599_o}),
    .q({open_n2008,\t/a/regfile/regfile$2$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1306 (
    .a({_al_u1302_o,_al_u1302_o}),
    .b({_al_u1303_o,_al_u1303_o}),
    .c({_al_u1304_o,_al_u1304_o}),
    .d({_al_u1305_o,_al_u1305_o}),
    .mi({open_n2021,\t/a/ID_rs2 [2]}),
    .fx({open_n2026,_al_u1306_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1311|t/a/regfile/reg0_b443  (
    .a({_al_u1306_o,_al_u1307_o}),
    .b({_al_u1308_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1310_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [27]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [27]}),
    .mi({open_n2030,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1311_o,_al_u1308_o}),
    .q({open_n2045,\t/a/regfile/regfile$13$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUT1("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .INIT_LUT0(16'b1011000000110000),
    .INIT_LUT1(16'b1111000001110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1317 (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .d({\t/a/regfile/regfile$31$ [27],\t/a/regfile/regfile$31$ [27]}),
    .mi({open_n2058,\t/a/regfile/regfile$30$ [27]}),
    .fx({open_n2063,_al_u1317_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1321|t/a/regfile/reg0_b955  (
    .a({_al_u1316_o,_al_u1317_o}),
    .b({_al_u1318_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1320_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [27]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [27]}),
    .mi({open_n2067,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1321_o,_al_u1318_o}),
    .q({open_n2082,\t/a/regfile/regfile$29$ [27]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1324|t/a/regfile/reg0_b986  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [26],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [26],\t/a/regfile/regfile$31$ [26]}),
    .e({open_n2083,\t/a/regfile/regfile$30$ [26]}),
    .mi({open_n2085,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1324_o,_al_u622_o}),
    .q({open_n2100,\t/a/regfile/regfile$30$ [26]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1332|t/a/regfile/reg0_b698  (
    .a({_al_u1327_o,_al_u1328_o}),
    .b({_al_u1329_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1331_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$20$ [26]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [26]}),
    .mi({open_n2102,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1332_o,_al_u1329_o}),
    .q({open_n2117,\t/a/regfile/regfile$21$ [26]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1336|t/a/regfile/reg0_b90  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [26],\t/a/regfile/regfile$3$ [26]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [26],\t/a/regfile/regfile$2$ [26]}),
    .mi({open_n2128,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1336_o,_al_u610_o}),
    .q({open_n2132,\t/a/regfile/regfile$2$ [26]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1337 (
    .a({_al_u1333_o,_al_u1333_o}),
    .b({_al_u1334_o,_al_u1334_o}),
    .c({_al_u1335_o,_al_u1335_o}),
    .d({_al_u1336_o,_al_u1336_o}),
    .mi({open_n2145,\t/a/ID_rs2 [2]}),
    .fx({open_n2150,_al_u1337_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1342|t/a/regfile/reg0_b442  (
    .a({_al_u1337_o,_al_u1338_o}),
    .b({_al_u1339_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1341_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [26]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [26]}),
    .mi({open_n2154,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1342_o,_al_u1339_o}),
    .q({open_n2169,\t/a/regfile/regfile$13$ [26]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1347|t/a/regfile/reg0_b89  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [25],\t/a/regfile/regfile$3$ [25]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [25],\t/a/regfile/regfile$2$ [25]}),
    .mi({open_n2180,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1347_o,_al_u631_o}),
    .q({open_n2184,\t/a/regfile/regfile$2$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1348 (
    .a({_al_u1344_o,_al_u1344_o}),
    .b({_al_u1345_o,_al_u1345_o}),
    .c({_al_u1346_o,_al_u1346_o}),
    .d({_al_u1347_o,_al_u1347_o}),
    .mi({open_n2197,\t/a/ID_rs2 [2]}),
    .fx({open_n2202,_al_u1348_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1353|t/a/regfile/reg0_b441  (
    .a({_al_u1348_o,_al_u1349_o}),
    .b({_al_u1350_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1352_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [25]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [25]}),
    .mi({open_n2206,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1353_o,_al_u1350_o}),
    .q({open_n2221,\t/a/regfile/regfile$13$ [25]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1011000000110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1111000001110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1359|t/a/regfile/reg0_b985  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$31$ [25],\t/a/regfile/regfile$31$ [25]}),
    .e({\t/a/regfile/regfile$30$ [25],\t/a/regfile/regfile$30$ [25]}),
    .mi({open_n2223,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1359_o,_al_u643_o}),
    .q({open_n2238,\t/a/regfile/regfile$30$ [25]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1363|t/a/regfile/reg0_b953  (
    .a({_al_u1358_o,_al_u1359_o}),
    .b({_al_u1360_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1362_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [25]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [25]}),
    .mi({open_n2240,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1363_o,_al_u1360_o}),
    .q({open_n2255,\t/a/regfile/regfile$29$ [25]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1365|t/a/regfile/reg0_b152  (
    .a({\t/a/ID_rs2 [0],_al_u2027_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$4$ [24],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [24],\t/a/reg_writedat [24]}),
    .mi({open_n2266,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1365_o,\t/a/aluin/sel1_b24/B9 }),
    .q({open_n2270,\t/a/regfile/regfile$4$ [24]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1368|t/a/regfile/reg0_b88  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [24],\t/a/regfile/regfile$3$ [24]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [24],\t/a/regfile/regfile$2$ [24]}),
    .mi({open_n2281,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1368_o,_al_u652_o}),
    .q({open_n2285,\t/a/regfile/regfile$2$ [24]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1374|t/a/regfile/reg0_b440  (
    .a({_al_u1369_o,_al_u1370_o}),
    .b({_al_u1371_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1373_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [24]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [24]}),
    .mi({open_n2287,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1374_o,_al_u1371_o}),
    .q({open_n2302,\t/a/regfile/regfile$13$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1379 (
    .a({_al_u1375_o,_al_u1375_o}),
    .b({_al_u1376_o,_al_u1376_o}),
    .c({_al_u1377_o,_al_u1377_o}),
    .d({_al_u1378_o,_al_u1378_o}),
    .mi({open_n2315,\t/a/ID_rs2 [2]}),
    .fx({open_n2320,_al_u1379_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1011000000110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1111000001110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1380|t/a/regfile/reg0_b984  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$31$ [24],\t/a/regfile/regfile$31$ [24]}),
    .e({\t/a/regfile/regfile$30$ [24],\t/a/regfile/regfile$30$ [24]}),
    .mi({open_n2324,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1380_o,_al_u664_o}),
    .q({open_n2339,\t/a/regfile/regfile$30$ [24]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1384|t/a/regfile/reg0_b952  (
    .a({_al_u1379_o,_al_u1380_o}),
    .b({_al_u1381_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1383_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [24]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [24]}),
    .mi({open_n2341,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1384_o,_al_u1381_o}),
    .q({open_n2356,\t/a/regfile/regfile$29$ [24]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1387|t/a/regfile/reg0_b983  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [23],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [23],\t/a/regfile/regfile$31$ [23]}),
    .e({open_n2357,\t/a/regfile/regfile$30$ [23]}),
    .mi({open_n2359,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1387_o,_al_u685_o}),
    .q({open_n2374,\t/a/regfile/regfile$30$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1390|_al_u1579  (
    .a({_al_u1386_o,_al_u1575_o}),
    .b({_al_u1387_o,_al_u1576_o}),
    .c({_al_u1388_o,_al_u1577_o}),
    .d({_al_u1389_o,_al_u1578_o}),
    .e({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .f({_al_u1390_o,_al_u1579_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1395|t/a/regfile/reg0_b695  (
    .a({_al_u1390_o,_al_u1391_o}),
    .b({_al_u1392_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1394_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$20$ [23]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [23]}),
    .mi({open_n2398,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1395_o,_al_u1392_o}),
    .q({open_n2413,\t/a/regfile/regfile$21$ [23]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1396|t/a/regfile/reg0_b151  (
    .a({\t/a/ID_rs2 [0],_al_u2030_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$4$ [23],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [23],\t/a/reg_writedat [23]}),
    .mi({open_n2417,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1396_o,\t/a/aluin/sel1_b23/B9 }),
    .q({open_n2432,\t/a/regfile/regfile$4$ [23]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1399|t/a/regfile/reg0_b87  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [23],\t/a/regfile/regfile$3$ [23]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [23],\t/a/regfile/regfile$2$ [23]}),
    .mi({open_n2443,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1399_o,_al_u673_o}),
    .q({open_n2447,\t/a/regfile/regfile$2$ [23]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1400 (
    .a({_al_u1396_o,_al_u1396_o}),
    .b({_al_u1397_o,_al_u1397_o}),
    .c({_al_u1398_o,_al_u1398_o}),
    .d({_al_u1399_o,_al_u1399_o}),
    .mi({open_n2460,\t/a/ID_rs2 [2]}),
    .fx({open_n2465,_al_u1400_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1405|t/a/regfile/reg0_b439  (
    .a({_al_u1400_o,_al_u1401_o}),
    .b({_al_u1402_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1404_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [23]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [23]}),
    .mi({open_n2469,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1405_o,_al_u1402_o}),
    .q({open_n2484,\t/a/regfile/regfile$13$ [23]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1407|t/a/regfile/reg0_b150  (
    .a({\t/a/ID_rs2 [0],_al_u2033_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$4$ [22],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [22],\t/a/reg_writedat [22]}),
    .mi({open_n2488,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1407_o,\t/a/aluin/sel1_b22/B9 }),
    .q({open_n2503,\t/a/regfile/regfile$4$ [22]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1410|t/a/regfile/reg0_b86  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [22],\t/a/regfile/regfile$3$ [22]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [22],\t/a/regfile/regfile$2$ [22]}),
    .mi({open_n2514,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1410_o,_al_u704_o}),
    .q({open_n2518,\t/a/regfile/regfile$2$ [22]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1416|t/a/regfile/reg0_b438  (
    .a({_al_u1411_o,_al_u1412_o}),
    .b({_al_u1413_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1415_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [22]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [22]}),
    .mi({open_n2520,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1416_o,_al_u1413_o}),
    .q({open_n2535,\t/a/regfile/regfile$13$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1011000000110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1111000001110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1422|_al_u1674  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .d({\t/a/regfile/regfile$31$ [22],\t/a/regfile/regfile$31$ [11]}),
    .e({\t/a/regfile/regfile$30$ [22],\t/a/regfile/regfile$30$ [11]}),
    .f({_al_u1422_o,_al_u1674_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1426|t/a/regfile/reg0_b950  (
    .a({_al_u1421_o,_al_u1422_o}),
    .b({_al_u1423_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1425_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [22]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [22]}),
    .mi({open_n2559,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1426_o,_al_u1423_o}),
    .q({open_n2574,\t/a/regfile/regfile$29$ [22]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1429|t/a/regfile/reg0_b981  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [21],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [21],\t/a/regfile/regfile$31$ [21]}),
    .e({open_n2575,\t/a/regfile/regfile$30$ [21]}),
    .mi({open_n2577,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1429_o,_al_u727_o}),
    .q({open_n2592,\t/a/regfile/regfile$30$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1432 (
    .a({_al_u1428_o,_al_u1428_o}),
    .b({_al_u1429_o,_al_u1429_o}),
    .c({_al_u1430_o,_al_u1430_o}),
    .d({_al_u1431_o,_al_u1431_o}),
    .mi({open_n2605,\t/a/ID_rs2 [2]}),
    .fx({open_n2610,_al_u1432_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1437|t/a/regfile/reg0_b693  (
    .a({_al_u1432_o,_al_u1433_o}),
    .b({_al_u1434_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1436_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$20$ [21]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [21]}),
    .mi({open_n2614,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1437_o,_al_u1434_o}),
    .q({open_n2629,\t/a/regfile/regfile$21$ [21]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1438|t/a/regfile/reg0_b149  (
    .a({\t/a/ID_rs2 [0],_al_u2036_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$4$ [21],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [21],\t/a/reg_writedat [21]}),
    .mi({open_n2640,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1438_o,\t/a/aluin/sel1_b21/B9 }),
    .q({open_n2644,\t/a/regfile/regfile$4$ [21]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1441|t/a/regfile/reg0_b85  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [21],\t/a/regfile/regfile$3$ [21]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [21],\t/a/regfile/regfile$2$ [21]}),
    .mi({open_n2655,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1441_o,_al_u715_o}),
    .q({open_n2659,\t/a/regfile/regfile$2$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1442 (
    .a({_al_u1438_o,_al_u1438_o}),
    .b({_al_u1439_o,_al_u1439_o}),
    .c({_al_u1440_o,_al_u1440_o}),
    .d({_al_u1441_o,_al_u1441_o}),
    .mi({open_n2672,\t/a/ID_rs2 [2]}),
    .fx({open_n2677,_al_u1442_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1447|t/a/regfile/reg0_b437  (
    .a({_al_u1442_o,_al_u1443_o}),
    .b({_al_u1444_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1446_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [21]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [21]}),
    .mi({open_n2681,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1447_o,_al_u1444_o}),
    .q({open_n2696,\t/a/regfile/regfile$13$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1449|_al_u1453  (
    .a({\t/a/ID_rs2 [0],_al_u1449_o}),
    .b({\t/a/ID_rs2 [1],_al_u1450_o}),
    .c({\t/a/regfile/regfile$4$ [20],_al_u1451_o}),
    .d({\t/a/regfile/regfile$5$ [20],_al_u1452_o}),
    .e({open_n2699,\t/a/ID_rs2 [2]}),
    .f({_al_u1449_o,_al_u1453_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1452|t/a/regfile/reg0_b84  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [20],\t/a/regfile/regfile$3$ [20]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [20],\t/a/regfile/regfile$2$ [20]}),
    .mi({open_n2730,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1452_o,_al_u746_o}),
    .q({open_n2734,\t/a/regfile/regfile$2$ [20]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1458|t/a/regfile/reg0_b436  (
    .a({_al_u1453_o,_al_u1454_o}),
    .b({_al_u1455_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1457_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [20]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [20]}),
    .mi({open_n2736,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1458_o,_al_u1455_o}),
    .q({open_n2751,\t/a/regfile/regfile$13$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1463|_al_u1464  (
    .a({_al_u1459_o,\t/a/ID_rs2 [0]}),
    .b({_al_u1460_o,\t/a/ID_rs2 [1]}),
    .c({_al_u1461_o,\t/a/ID_rs2 [2]}),
    .d({_al_u1462_o,\t/a/regfile/regfile$31$ [20]}),
    .e({\t/a/ID_rs2 [2],\t/a/regfile/regfile$30$ [20]}),
    .f({_al_u1463_o,_al_u1464_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1468|t/a/regfile/reg0_b948  (
    .a({_al_u1463_o,_al_u1464_o}),
    .b({_al_u1465_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1467_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [20]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [20]}),
    .mi({open_n2775,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1468_o,_al_u1465_o}),
    .q({open_n2790,\t/a/regfile/regfile$29$ [20]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(C*~(D*~A*~(~0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~(C*~(D*~A*~(~1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001111100001111),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0101111100001111),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1470|t/a/regfile/reg0_b161  (
    .a({\t/a/ID_rs2 [0],_al_u2072_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$4$ [1],_al_u2073_o}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [1],\t/a/aluin/n10_lutinv }),
    .e({open_n2791,\t/a/reg_writedat [1]}),
    .mi({open_n2793,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u1470_o,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .q({open_n2808,\t/a/regfile/regfile$5$ [1]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1471|_al_u1474  (
    .a({\t/a/ID_rs2 [0],_al_u1470_o}),
    .b({\t/a/ID_rs2 [1],_al_u1471_o}),
    .c({\t/a/regfile/regfile$6$ [1],_al_u1472_o}),
    .d({\t/a/regfile/regfile$7$ [1],_al_u1473_o}),
    .e({open_n2811,\t/a/ID_rs2 [2]}),
    .f({_al_u1471_o,_al_u1474_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1479|t/a/regfile/reg0_b417  (
    .a({_al_u1474_o,_al_u1475_o}),
    .b({_al_u1476_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1478_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [1]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [1]}),
    .mi({open_n2833,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u1479_o,_al_u1476_o}),
    .q({open_n2848,\t/a/regfile/regfile$13$ [1]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1484 (
    .a({_al_u1480_o,_al_u1480_o}),
    .b({_al_u1481_o,_al_u1481_o}),
    .c({_al_u1482_o,_al_u1482_o}),
    .d({_al_u1483_o,_al_u1483_o}),
    .mi({open_n2861,\t/a/ID_rs2 [2]}),
    .fx({open_n2866,_al_u1484_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1489|t/a/regfile/reg0_b929  (
    .a({_al_u1484_o,_al_u1485_o}),
    .b({_al_u1486_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1488_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [1]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [1]}),
    .mi({open_n2870,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u1489_o,_al_u1486_o}),
    .q({open_n2885,\t/a/regfile/regfile$29$ [1]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1491|t/a/regfile/reg0_b147  (
    .a({\t/a/ID_rs2 [0],_al_u2042_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$4$ [19],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [19],\t/a/reg_writedat [19]}),
    .mi({open_n2889,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1491_o,\t/a/aluin/sel1_b19/B9 }),
    .q({open_n2904,\t/a/regfile/regfile$4$ [19]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1494|t/a/regfile/reg0_b83  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [19],\t/a/regfile/regfile$3$ [19]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [19],\t/a/regfile/regfile$2$ [19]}),
    .mi({open_n2915,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1494_o,_al_u778_o}),
    .q({open_n2919,\t/a/regfile/regfile$2$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1495 (
    .a({_al_u1491_o,_al_u1491_o}),
    .b({_al_u1492_o,_al_u1492_o}),
    .c({_al_u1493_o,_al_u1493_o}),
    .d({_al_u1494_o,_al_u1494_o}),
    .mi({open_n2932,\t/a/ID_rs2 [2]}),
    .fx({open_n2937,_al_u1495_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1500|t/a/regfile/reg0_b435  (
    .a({_al_u1495_o,_al_u1496_o}),
    .b({_al_u1497_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1499_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [19]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [19]}),
    .mi({open_n2941,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1500_o,_al_u1497_o}),
    .q({open_n2956,\t/a/regfile/regfile$13$ [19]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1011000000110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1111000001110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1506|t/a/regfile/reg0_b979  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$31$ [19],\t/a/regfile/regfile$31$ [19]}),
    .e({\t/a/regfile/regfile$30$ [19],\t/a/regfile/regfile$30$ [19]}),
    .mi({open_n2958,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1506_o,_al_u790_o}),
    .q({open_n2973,\t/a/regfile/regfile$30$ [19]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1510|t/a/regfile/reg0_b947  (
    .a({_al_u1505_o,_al_u1506_o}),
    .b({_al_u1507_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1509_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [19]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [19]}),
    .mi({open_n2975,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1510_o,_al_u1507_o}),
    .q({open_n2990,\t/a/regfile/regfile$29$ [19]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1512|t/a/regfile/reg0_b146  (
    .a({\t/a/ID_rs2 [0],_al_u2045_o}),
    .b({\t/a/ID_rs2 [1],\t/a/alu_B_select [1]}),
    .c({\t/a/regfile/regfile$4$ [18],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [18],\t/a/reg_writedat [18]}),
    .mi({open_n2994,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1512_o,\t/a/aluin/sel1_b18/B9 }),
    .q({open_n3009,\t/a/regfile/regfile$4$ [18]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1515|t/a/regfile/reg0_b82  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [18],\t/a/regfile/regfile$3$ [18]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [18],\t/a/regfile/regfile$2$ [18]}),
    .mi({open_n3020,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1515_o,_al_u809_o}),
    .q({open_n3024,\t/a/regfile/regfile$2$ [18]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1521|t/a/regfile/reg0_b434  (
    .a({_al_u1516_o,_al_u1517_o}),
    .b({_al_u1518_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1520_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [18]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [18]}),
    .mi({open_n3026,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1521_o,_al_u1518_o}),
    .q({open_n3041,\t/a/regfile/regfile$13$ [18]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1526|_al_u1527  (
    .a({_al_u1522_o,\t/a/ID_rs2 [0]}),
    .b({_al_u1523_o,\t/a/ID_rs2 [1]}),
    .c({_al_u1524_o,\t/a/ID_rs2 [2]}),
    .d({_al_u1525_o,\t/a/regfile/regfile$31$ [18]}),
    .e({\t/a/ID_rs2 [2],\t/a/regfile/regfile$30$ [18]}),
    .f({_al_u1526_o,_al_u1527_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1531|t/a/regfile/reg0_b946  (
    .a({_al_u1526_o,_al_u1527_o}),
    .b({_al_u1528_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1530_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [18]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [18]}),
    .mi({open_n3065,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1531_o,_al_u1528_o}),
    .q({open_n3080,\t/a/regfile/regfile$29$ [18]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1534|t/a/regfile/reg0_b977  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [17],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [17],\t/a/regfile/regfile$31$ [17]}),
    .e({open_n3081,\t/a/regfile/regfile$30$ [17]}),
    .mi({open_n3083,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1534_o,_al_u832_o}),
    .q({open_n3098,\t/a/regfile/regfile$30$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1537 (
    .a({_al_u1533_o,_al_u1533_o}),
    .b({_al_u1534_o,_al_u1534_o}),
    .c({_al_u1535_o,_al_u1535_o}),
    .d({_al_u1536_o,_al_u1536_o}),
    .mi({open_n3111,\t/a/ID_rs2 [2]}),
    .fx({open_n3116,_al_u1537_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1542|t/a/regfile/reg0_b689  (
    .a({_al_u1537_o,_al_u1538_o}),
    .b({_al_u1539_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1541_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$20$ [17]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [17]}),
    .mi({open_n3120,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1542_o,_al_u1539_o}),
    .q({open_n3135,\t/a/regfile/regfile$21$ [17]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1543|t/a/regfile/reg0_b945  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$4$ [17],\t/a/regfile/regfile$28$ [17]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [17],\t/a/regfile/regfile$29$ [17]}),
    .mi({open_n3146,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1543_o,_al_u1533_o}),
    .q({open_n3150,\t/a/regfile/regfile$29$ [17]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1545|t/a/regfile/reg0_b49  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$0$ [17],\t/a/regfile/regfile$0$ [17]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [17],\t/a/regfile/regfile$1$ [17]}),
    .mi({open_n3161,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1545_o,_al_u819_o}),
    .q({open_n3165,\t/a/regfile/regfile$1$ [17]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1546|t/a/regfile/reg0_b81  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [17],\t/a/regfile/regfile$3$ [17]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [17],\t/a/regfile/regfile$2$ [17]}),
    .mi({open_n3176,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1546_o,_al_u820_o}),
    .q({open_n3180,\t/a/regfile/regfile$2$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1547 (
    .a({_al_u1543_o,_al_u1543_o}),
    .b({_al_u1544_o,_al_u1544_o}),
    .c({_al_u1545_o,_al_u1545_o}),
    .d({_al_u1546_o,_al_u1546_o}),
    .mi({open_n3193,\t/a/ID_rs2 [2]}),
    .fx({open_n3198,_al_u1547_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1552|t/a/regfile/reg0_b433  (
    .a({_al_u1547_o,_al_u1548_o}),
    .b({_al_u1549_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1551_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [17]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [17]}),
    .mi({open_n3202,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1552_o,_al_u1549_o}),
    .q({open_n3217,\t/a/regfile/regfile$13$ [17]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1554|t/a/regfile/reg0_b240  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$4$ [16],\t/a/regfile/regfile$6$ [16]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [16],\t/a/regfile/regfile$7$ [16]}),
    .mi({open_n3228,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1554_o,_al_u1555_o}),
    .q({open_n3232,\t/a/regfile/regfile$7$ [16]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1556|t/a/regfile/reg0_b48  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$0$ [16],\t/a/regfile/regfile$0$ [16]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [16],\t/a/regfile/regfile$1$ [16]}),
    .mi({open_n3243,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1556_o,_al_u850_o}),
    .q({open_n3247,\t/a/regfile/regfile$1$ [16]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1557|t/a/regfile/reg0_b80  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [16],\t/a/regfile/regfile$3$ [16]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [16],\t/a/regfile/regfile$2$ [16]}),
    .mi({open_n3258,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1557_o,_al_u851_o}),
    .q({open_n3262,\t/a/regfile/regfile$2$ [16]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1563|t/a/regfile/reg0_b432  (
    .a({_al_u1558_o,_al_u1559_o}),
    .b({_al_u1560_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1562_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [16]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [16]}),
    .mi({open_n3264,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1563_o,_al_u1560_o}),
    .q({open_n3279,\t/a/regfile/regfile$13$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1568|_al_u1610  (
    .a({_al_u1564_o,_al_u1606_o}),
    .b({_al_u1565_o,_al_u1607_o}),
    .c({_al_u1566_o,_al_u1608_o}),
    .d({_al_u1567_o,_al_u1609_o}),
    .e({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .f({_al_u1568_o,_al_u1610_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUT1("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .INIT_LUT0(16'b1011000000110000),
    .INIT_LUT1(16'b1111000001110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1569 (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .d({\t/a/regfile/regfile$31$ [16],\t/a/regfile/regfile$31$ [16]}),
    .mi({open_n3314,\t/a/regfile/regfile$30$ [16]}),
    .fx({open_n3319,_al_u1569_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1573|t/a/regfile/reg0_b944  (
    .a({_al_u1568_o,_al_u1569_o}),
    .b({_al_u1570_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1572_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [16]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [16]}),
    .mi({open_n3323,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1573_o,_al_u1570_o}),
    .q({open_n3338,\t/a/regfile/regfile$29$ [16]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1576|t/a/regfile/reg0_b975  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [15],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [15],\t/a/regfile/regfile$31$ [15]}),
    .e({open_n3339,\t/a/regfile/regfile$30$ [15]}),
    .mi({open_n3341,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1576_o,_al_u874_o}),
    .q({open_n3356,\t/a/regfile/regfile$30$ [15]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1584|t/a/regfile/reg0_b687  (
    .a({_al_u1579_o,_al_u1580_o}),
    .b({_al_u1581_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1583_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$20$ [15]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [15]}),
    .mi({open_n3358,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1584_o,_al_u1581_o}),
    .q({open_n3373,\t/a/regfile/regfile$21$ [15]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1585|t/a/regfile/reg0_b175  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$4$ [15],\t/a/regfile/regfile$4$ [15]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [15],\t/a/regfile/regfile$5$ [15]}),
    .mi({open_n3384,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1585_o,_al_u859_o}),
    .q({open_n3388,\t/a/regfile/regfile$5$ [15]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1587|t/a/regfile/reg0_b47  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$0$ [15],\t/a/regfile/regfile$0$ [15]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [15],\t/a/regfile/regfile$1$ [15]}),
    .mi({open_n3399,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1587_o,_al_u861_o}),
    .q({open_n3403,\t/a/regfile/regfile$1$ [15]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1588|t/a/regfile/reg0_b79  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [15],\t/a/regfile/regfile$3$ [15]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [15],\t/a/regfile/regfile$2$ [15]}),
    .mi({open_n3414,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1588_o,_al_u862_o}),
    .q({open_n3418,\t/a/regfile/regfile$2$ [15]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1589 (
    .a({_al_u1585_o,_al_u1585_o}),
    .b({_al_u1586_o,_al_u1586_o}),
    .c({_al_u1587_o,_al_u1587_o}),
    .d({_al_u1588_o,_al_u1588_o}),
    .mi({open_n3431,\t/a/ID_rs2 [2]}),
    .fx({open_n3436,_al_u1589_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1594|t/a/regfile/reg0_b431  (
    .a({_al_u1589_o,_al_u1590_o}),
    .b({_al_u1591_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1593_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [15]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [15]}),
    .mi({open_n3440,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1594_o,_al_u1591_o}),
    .q({open_n3455,\t/a/regfile/regfile$13$ [15]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1596|t/a/regfile/reg0_b174  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$4$ [14],\t/a/regfile/regfile$4$ [14]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [14],\t/a/regfile/regfile$5$ [14]}),
    .mi({open_n3466,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1596_o,_al_u880_o}),
    .q({open_n3470,\t/a/regfile/regfile$5$ [14]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1598|_al_u1516  (
    .a({\t/a/ID_rs2 [0],_al_u1512_o}),
    .b({\t/a/ID_rs2 [1],_al_u1513_o}),
    .c({\t/a/regfile/regfile$0$ [14],_al_u1514_o}),
    .d({\t/a/regfile/regfile$1$ [14],_al_u1515_o}),
    .e({open_n3473,\t/a/ID_rs2 [2]}),
    .f({_al_u1598_o,_al_u1516_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1599|t/a/regfile/reg0_b78  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [14],\t/a/regfile/regfile$3$ [14]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [14],\t/a/regfile/regfile$2$ [14]}),
    .mi({open_n3504,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1599_o,_al_u883_o}),
    .q({open_n3508,\t/a/regfile/regfile$2$ [14]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1600 (
    .a({_al_u1596_o,_al_u1596_o}),
    .b({_al_u1597_o,_al_u1597_o}),
    .c({_al_u1598_o,_al_u1598_o}),
    .d({_al_u1599_o,_al_u1599_o}),
    .mi({open_n3521,\t/a/ID_rs2 [2]}),
    .fx({open_n3526,_al_u1600_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1605|t/a/regfile/reg0_b430  (
    .a({_al_u1600_o,_al_u1601_o}),
    .b({_al_u1602_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1604_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [14]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [14]}),
    .mi({open_n3530,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1605_o,_al_u1602_o}),
    .q({open_n3545,\t/a/regfile/regfile$13$ [14]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1011000000110000),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1111000001110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1611|t/a/regfile/reg0_b974  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$31$ [14],\t/a/regfile/regfile$31$ [14]}),
    .e({\t/a/regfile/regfile$30$ [14],\t/a/regfile/regfile$30$ [14]}),
    .mi({open_n3547,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1611_o,_al_u895_o}),
    .q({open_n3562,\t/a/regfile/regfile$30$ [14]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1615|t/a/regfile/reg0_b942  (
    .a({_al_u1610_o,_al_u1611_o}),
    .b({_al_u1612_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1614_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [14]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [14]}),
    .mi({open_n3564,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1615_o,_al_u1612_o}),
    .q({open_n3579,\t/a/regfile/regfile$29$ [14]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1617|t/a/regfile/reg0_b173  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$4$ [13],\t/a/regfile/regfile$4$ [13]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [13],\t/a/regfile/regfile$5$ [13]}),
    .mi({open_n3590,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1617_o,_al_u911_o}),
    .q({open_n3594,\t/a/regfile/regfile$5$ [13]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1619|_al_u1621  (
    .a({\t/a/ID_rs2 [0],_al_u1617_o}),
    .b({\t/a/ID_rs2 [1],_al_u1618_o}),
    .c({\t/a/regfile/regfile$0$ [13],_al_u1619_o}),
    .d({\t/a/regfile/regfile$1$ [13],_al_u1620_o}),
    .e({open_n3597,\t/a/ID_rs2 [2]}),
    .f({_al_u1619_o,_al_u1621_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1620|t/a/regfile/reg0_b77  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [13],\t/a/regfile/regfile$3$ [13]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [13],\t/a/regfile/regfile$2$ [13]}),
    .mi({open_n3628,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1620_o,_al_u914_o}),
    .q({open_n3632,\t/a/regfile/regfile$2$ [13]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1626|t/a/regfile/reg0_b429  (
    .a({_al_u1621_o,_al_u1622_o}),
    .b({_al_u1623_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1625_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [13]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [13]}),
    .mi({open_n3634,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1626_o,_al_u1623_o}),
    .q({open_n3649,\t/a/regfile/regfile$13$ [13]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1631 (
    .a({_al_u1627_o,_al_u1627_o}),
    .b({_al_u1628_o,_al_u1628_o}),
    .c({_al_u1629_o,_al_u1629_o}),
    .d({_al_u1630_o,_al_u1630_o}),
    .mi({open_n3662,\t/a/ID_rs2 [2]}),
    .fx({open_n3667,_al_u1631_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUT1("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    .INIT_LUT0(16'b1011000000110000),
    .INIT_LUT1(16'b1111000001110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1632 (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .d({\t/a/regfile/regfile$31$ [13],\t/a/regfile/regfile$31$ [13]}),
    .mi({open_n3682,\t/a/regfile/regfile$30$ [13]}),
    .fx({open_n3687,_al_u1632_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1636|t/a/regfile/reg0_b941  (
    .a({_al_u1631_o,_al_u1632_o}),
    .b({_al_u1633_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1635_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [13]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [13]}),
    .mi({open_n3691,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1636_o,_al_u1633_o}),
    .q({open_n3706,\t/a/regfile/regfile$29$ [13]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1639|t/a/regfile/reg0_b972  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [12],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [12],\t/a/regfile/regfile$31$ [12]}),
    .e({open_n3707,\t/a/regfile/regfile$30$ [12]}),
    .mi({open_n3709,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1639_o,_al_u937_o}),
    .q({open_n3724,\t/a/regfile/regfile$30$ [12]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1642 (
    .a({_al_u1638_o,_al_u1638_o}),
    .b({_al_u1639_o,_al_u1639_o}),
    .c({_al_u1640_o,_al_u1640_o}),
    .d({_al_u1641_o,_al_u1641_o}),
    .mi({open_n3737,\t/a/ID_rs2 [2]}),
    .fx({open_n3742,_al_u1642_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1647|t/a/regfile/reg0_b684  (
    .a({_al_u1642_o,_al_u1643_o}),
    .b({_al_u1644_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1646_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$20$ [12]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [12]}),
    .mi({open_n3746,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1647_o,_al_u1644_o}),
    .q({open_n3761,\t/a/regfile/regfile$21$ [12]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1648|t/a/regfile/reg0_b172  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$4$ [12],\t/a/regfile/regfile$4$ [12]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [12],\t/a/regfile/regfile$5$ [12]}),
    .mi({open_n3772,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1648_o,_al_u922_o}),
    .q({open_n3776,\t/a/regfile/regfile$5$ [12]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1650|_al_u1652  (
    .a({\t/a/ID_rs2 [0],_al_u1648_o}),
    .b({\t/a/ID_rs2 [1],_al_u1649_o}),
    .c({\t/a/regfile/regfile$0$ [12],_al_u1650_o}),
    .d({\t/a/regfile/regfile$1$ [12],_al_u1651_o}),
    .e({open_n3779,\t/a/ID_rs2 [2]}),
    .f({_al_u1650_o,_al_u1652_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1651|t/a/regfile/reg0_b76  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [12],\t/a/regfile/regfile$3$ [12]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [12],\t/a/regfile/regfile$2$ [12]}),
    .mi({open_n3810,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1651_o,_al_u925_o}),
    .q({open_n3814,\t/a/regfile/regfile$2$ [12]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1657|t/a/regfile/reg0_b428  (
    .a({_al_u1652_o,_al_u1653_o}),
    .b({_al_u1654_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1656_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [12]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [12]}),
    .mi({open_n3816,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1657_o,_al_u1654_o}),
    .q({open_n3831,\t/a/regfile/regfile$13$ [12]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1659|t/a/regfile/reg0_b171  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$4$ [11],\t/a/regfile/regfile$4$ [11]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [11],\t/a/regfile/regfile$5$ [11]}),
    .mi({open_n3842,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u1659_o,_al_u953_o}),
    .q({open_n3846,\t/a/regfile/regfile$5$ [11]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1661|_al_u1663  (
    .a({\t/a/ID_rs2 [0],_al_u1659_o}),
    .b({\t/a/ID_rs2 [1],_al_u1660_o}),
    .c({\t/a/regfile/regfile$0$ [11],_al_u1661_o}),
    .d({\t/a/regfile/regfile$1$ [11],_al_u1662_o}),
    .e({open_n3849,\t/a/ID_rs2 [2]}),
    .f({_al_u1661_o,_al_u1663_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1662|t/a/regfile/reg0_b75  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [11],\t/a/regfile/regfile$3$ [11]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [11],\t/a/regfile/regfile$2$ [11]}),
    .mi({open_n3880,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u1662_o,_al_u956_o}),
    .q({open_n3884,\t/a/regfile/regfile$2$ [11]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1668|t/a/regfile/reg0_b427  (
    .a({_al_u1663_o,_al_u1664_o}),
    .b({_al_u1665_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1667_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [11]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [11]}),
    .mi({open_n3886,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u1668_o,_al_u1665_o}),
    .q({open_n3901,\t/a/regfile/regfile$13$ [11]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1673 (
    .a({_al_u1669_o,_al_u1669_o}),
    .b({_al_u1670_o,_al_u1670_o}),
    .c({_al_u1671_o,_al_u1671_o}),
    .d({_al_u1672_o,_al_u1672_o}),
    .mi({open_n3914,\t/a/ID_rs2 [2]}),
    .fx({open_n3919,_al_u1673_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1678|t/a/regfile/reg0_b939  (
    .a({_al_u1673_o,_al_u1674_o}),
    .b({_al_u1675_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1677_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$28$ [11]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$29$ [11]}),
    .mi({open_n3923,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u1678_o,_al_u1675_o}),
    .q({open_n3938,\t/a/regfile/regfile$29$ [11]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b0000100001001100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b0000100001001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1681|t/a/regfile/reg0_b970  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [10],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [10],\t/a/regfile/regfile$31$ [10]}),
    .e({open_n3939,\t/a/regfile/regfile$30$ [10]}),
    .mi({open_n3941,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1681_o,_al_u979_o}),
    .q({open_n3956,\t/a/regfile/regfile$30$ [10]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1684 (
    .a({_al_u1680_o,_al_u1680_o}),
    .b({_al_u1681_o,_al_u1681_o}),
    .c({_al_u1682_o,_al_u1682_o}),
    .d({_al_u1683_o,_al_u1683_o}),
    .mi({open_n3969,\t/a/ID_rs2 [2]}),
    .fx({open_n3974,_al_u1684_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1689|t/a/regfile/reg0_b682  (
    .a({_al_u1684_o,_al_u1685_o}),
    .b({_al_u1686_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1688_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$20$ [10]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$21$ [10]}),
    .mi({open_n3978,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1689_o,_al_u1686_o}),
    .q({open_n3993,\t/a/regfile/regfile$21$ [10]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1690|t/a/regfile/reg0_b170  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$4$ [10],\t/a/regfile/regfile$4$ [10]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [10],\t/a/regfile/regfile$5$ [10]}),
    .mi({open_n4004,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1690_o,_al_u964_o}),
    .q({open_n4008,\t/a/regfile/regfile$5$ [10]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1692|_al_u1694  (
    .a({\t/a/ID_rs2 [0],_al_u1690_o}),
    .b({\t/a/ID_rs2 [1],_al_u1691_o}),
    .c({\t/a/regfile/regfile$0$ [10],_al_u1692_o}),
    .d({\t/a/regfile/regfile$1$ [10],_al_u1693_o}),
    .e({open_n4011,\t/a/ID_rs2 [2]}),
    .f({_al_u1692_o,_al_u1694_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1693|t/a/regfile/reg0_b74  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$3$ [10],\t/a/regfile/regfile$3$ [10]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$2$ [10],\t/a/regfile/regfile$2$ [10]}),
    .mi({open_n4042,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1693_o,_al_u967_o}),
    .q({open_n4046,\t/a/regfile/regfile$2$ [10]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1699|t/a/regfile/reg0_b426  (
    .a({_al_u1694_o,_al_u1695_o}),
    .b({_al_u1696_o,\t/a/ID_rs2 [0]}),
    .c({_al_u1698_o,\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs2 [3],\t/a/regfile/regfile$12$ [10]}),
    .e({\t/a/ID_rs2 [4],\t/a/regfile/regfile$13$ [10]}),
    .mi({open_n4048,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1699_o,_al_u1696_o}),
    .q({open_n4063,\t/a/regfile/regfile$13$ [10]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*~C*B*A)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~1*D*~C*B*A)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1701|t/a/regfile/reg0_b160  (
    .a({\t/a/ID_rs2 [0],_al_u254_o}),
    .b({\t/a/ID_rs2 [1],\t/a/WB_rd [0]}),
    .c({\t/a/regfile/regfile$4$ [0],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [0],\t/a/WB_rd [2]}),
    .e({open_n4064,\t/a/WB_rd [3]}),
    .mi({open_n4066,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1701_o,\t/a/regfile/mux39_b160_sel_is_3_o }),
    .q({open_n4081,\t/a/regfile/regfile$5$ [0]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*C*B*A)"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~1*D*C*B*A)"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1702|t/a/regfile/reg0_b224  (
    .a({\t/a/ID_rs2 [0],_al_u254_o}),
    .b({\t/a/ID_rs2 [1],\t/a/WB_rd [0]}),
    .c({\t/a/regfile/regfile$6$ [0],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [0],\t/a/WB_rd [2]}),
    .e({open_n4082,\t/a/WB_rd [3]}),
    .mi({open_n4084,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1702_o,\t/a/regfile/mux39_b224_sel_is_3_o }),
    .q({open_n4099,\t/a/regfile/regfile$7$ [0]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*B*A)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~1*~D*~C*B*A)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1703|t/a/regfile/reg0_b32  (
    .a({\t/a/ID_rs2 [0],_al_u254_o}),
    .b({\t/a/ID_rs2 [1],\t/a/WB_rd [0]}),
    .c({\t/a/regfile/regfile$0$ [0],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [0],\t/a/WB_rd [2]}),
    .e({open_n4100,\t/a/WB_rd [3]}),
    .mi({open_n4102,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1703_o,\t/a/regfile/mux39_b32_sel_is_3_o }),
    .q({open_n4117,\t/a/regfile/regfile$1$ [0]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*C*~B*A)"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~1*~D*C*~B*A)"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1704|t/a/regfile/reg0_b64  (
    .a({\t/a/ID_rs2 [0],_al_u254_o}),
    .b({\t/a/ID_rs2 [1],\t/a/WB_rd [0]}),
    .c({\t/a/regfile/regfile$2$ [0],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$3$ [0],\t/a/WB_rd [2]}),
    .e({open_n4118,\t/a/WB_rd [3]}),
    .mi({open_n4120,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1704_o,\t/a/regfile/mux39_b64_sel_is_3_o }),
    .q({open_n4135,\t/a/regfile/regfile$2$ [0]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*B*A)"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(1*D*~C*B*A)"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1707|t/a/regfile/reg0_b416  (
    .a({_al_u1706_o,_al_u254_o}),
    .b({\t/a/ID_rs2 [0],\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$12$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$13$ [0],\t/a/WB_rd [3]}),
    .mi({open_n4137,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1707_o,\t/a/regfile/mux39_b416_sel_is_3_o }),
    .q({open_n4152,\t/a/regfile/regfile$13$ [0]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUT1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUT0(16'b0000011100000011),
    .INIT_LUT1(16'b0000111100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1708 (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .d({\t/a/regfile/regfile$10$ [0],\t/a/regfile/regfile$10$ [0]}),
    .mi({open_n4165,\t/a/regfile/regfile$11$ [0]}),
    .fx({open_n4170,_al_u1708_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUT1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .INIT_LUT0(16'b1010001010100000),
    .INIT_LUT1(16'b1010101010101000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1709 (
    .a({_al_u1708_o,_al_u1708_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .d({\t/a/regfile/regfile$8$ [0],\t/a/regfile/regfile$8$ [0]}),
    .mi({open_n4185,\t/a/regfile/regfile$9$ [0]}),
    .fx({open_n4190,_al_u1709_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1710|_al_u1705  (
    .a({_al_u1705_o,_al_u1701_o}),
    .b({_al_u1707_o,_al_u1702_o}),
    .c({_al_u1709_o,_al_u1703_o}),
    .d({\t/a/ID_rs2 [3],_al_u1704_o}),
    .e({\t/a/ID_rs2 [4],\t/a/ID_rs2 [2]}),
    .f({_al_u1710_o,_al_u1705_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*~C*B*A)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~1*D*~C*B*A)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1711|t/a/regfile/reg0_b672  (
    .a({\t/a/ID_rs2 [0],_al_u256_o}),
    .b({\t/a/ID_rs2 [1],\t/a/WB_rd [0]}),
    .c({\t/a/regfile/regfile$20$ [0],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [0],\t/a/WB_rd [2]}),
    .e({open_n4215,\t/a/WB_rd [3]}),
    .mi({open_n4217,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1711_o,\t/a/regfile/mux39_b672_sel_is_3_o }),
    .q({open_n4232,\t/a/regfile/regfile$21$ [0]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1715 (
    .a({_al_u1711_o,_al_u1711_o}),
    .b({_al_u1712_o,_al_u1712_o}),
    .c({_al_u1713_o,_al_u1713_o}),
    .d({_al_u1714_o,_al_u1714_o}),
    .mi({open_n4245,\t/a/ID_rs2 [2]}),
    .fx({open_n4250,_al_u1715_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUT1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUT0(16'b0111000000110000),
    .INIT_LUT1(16'b1111000010110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1716 (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .d({\t/a/regfile/regfile$30$ [0],\t/a/regfile/regfile$30$ [0]}),
    .mi({open_n4265,\t/a/regfile/regfile$31$ [0]}),
    .fx({open_n4270,_al_u1716_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*~B*A)"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(1*D*~C*~B*A)"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1717|t/a/regfile/reg0_b896  (
    .a({_al_u1716_o,_al_u256_o}),
    .b({\t/a/ID_rs2 [0],\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$28$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$29$ [0],\t/a/WB_rd [3]}),
    .mi({open_n4274,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1717_o,\t/a/regfile/mux39_b896_sel_is_3_o }),
    .q({open_n4289,\t/a/regfile/regfile$28$ [0]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUT1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .INIT_LUT0(16'b1010001010100000),
    .INIT_LUT1(16'b1010101010101000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1719 (
    .a({_al_u1718_o,_al_u1718_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .d({\t/a/regfile/regfile$24$ [0],\t/a/regfile/regfile$24$ [0]}),
    .mi({open_n4302,\t/a/regfile/regfile$25$ [0]}),
    .fx({open_n4307,_al_u1719_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1722|_al_u1723  (
    .a({\t/a/MEM_rd [1],_al_u1722_o}),
    .b({\t/a/MEM_rd [2],\t/a/MEM_rd [3]}),
    .c({\t/a/ID_rs2 [1],\t/a/MEM_rd [4]}),
    .d({\t/a/ID_rs2 [2],\t/a/ID_rs2 [3]}),
    .e({open_n4312,\t/a/ID_rs2 [4]}),
    .f({_al_u1722_o,_al_u1723_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1726|_al_u1725  (
    .a({open_n4333,_al_u1724_o}),
    .b({open_n4334,\t/a/MEM_rd [0]}),
    .c({_al_u1725_o,\t/a/MEM_rd [1]}),
    .d({_al_u1723_o,\t/a/ID_rs2 [0]}),
    .e({open_n4337,\t/a/ID_rs2 [1]}),
    .f({\t/a/risk_jump/n42_lutinv ,_al_u1725_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1730|_al_u348  (
    .a({\t/a/MEM_rd [1],_al_u344_o}),
    .b({\t/a/MEM_rd [3],_al_u345_o}),
    .c({\t/a/ID_rs1 [1],_al_u346_o}),
    .d({\t/a/ID_rs1 [3],_al_u347_o}),
    .e({open_n4360,\t/a/ID_rs1 [2]}),
    .f({_al_u1730_o,_al_u348_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1731|_al_u1728  (
    .a({_al_u1728_o,_al_u1727_o}),
    .b({_al_u1729_o,\t/a/MEM_rd [0]}),
    .c({_al_u1730_o,\t/a/MEM_rd [2]}),
    .d({\t/a/MEM_rd [4],\t/a/ID_rs1 [0]}),
    .e({\t/a/ID_rs1 [4],\t/a/ID_rs1 [2]}),
    .f({\t/a/risk_jump/n24_lutinv ,_al_u1728_o}));
  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(~D*~C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1732|t/a/mem_wb/reg1_b5  (
    .a({_al_u251_o,_al_u251_o}),
    .b({_al_u252_o,_al_u252_o}),
    .c({\t/a/MEM_op [5],\t/a/MEM_op [5]}),
    .ce(\t/a/ex_mem/n0 ),
    .clk(clock_pad),
    .d({\t/a/MEM_op [6],\t/a/MEM_op [6]}),
    .mi({open_n4413,\t/a/MEM_op [5]}),
    .f({\t/busarbitration/mux5_b0_sel_is_3_o ,memwrite_cs}),
    .q({open_n4418,\t/a/WB_op [5]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b0000001110101010),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1734|_al_u1720  (
    .a({\t/a/EX_rd [0],_al_u1715_o}),
    .b({\t/a/EX_rd [1],_al_u1717_o}),
    .c({\t/a/ID_rs2 [0],_al_u1719_o}),
    .d({\t/a/ID_rs2 [1],\t/a/ID_rs2 [3]}),
    .e({open_n4421,\t/a/ID_rs2 [4]}),
    .f({_al_u1734_o,_al_u1720_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(0@C)*~(D@B))"),
    //.LUT1("(A*~(1@C)*~(D@B))"),
    .INIT_LUT0(16'b0000100000000010),
    .INIT_LUT1(16'b1000000000100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1735 (
    .a({_al_u1734_o,_al_u1734_o}),
    .b({\t/a/EX_rd [3],\t/a/EX_rd [3]}),
    .c({\t/a/EX_rd [4],\t/a/EX_rd [4]}),
    .d({\t/a/ID_rs2 [3],\t/a/ID_rs2 [3]}),
    .mi({open_n4454,\t/a/ID_rs2 [4]}),
    .fx({open_n4459,_al_u1735_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0@C)*~(D*~B))"),
    //.LUT1("(~A*~(1@C)*~(D*~B))"),
    .INIT_LUT0(16'b0000010000000101),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1737 (
    .a({_al_u1736_o,_al_u1736_o}),
    .b({\t/a/EX_rd [0],\t/a/EX_rd [0]}),
    .c({\t/a/EX_rd [2],\t/a/EX_rd [2]}),
    .d({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .mi({open_n4474,\t/a/ID_rs2 [2]}),
    .fx({open_n4479,_al_u1737_o}));
  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~B*~(D*A)))"),
    //.LUT1("(~C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110000011000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1740|t/a/ex_mem/reg2_b4  (
    .a({open_n4482,_al_u1984_o}),
    .b({\t/a/EX_op [3],\t/a/aluin/n10_lutinv }),
    .c({\t/a/EX_op [4],\t/a/EX_fun3 [1]}),
    .clk(clock_pad),
    .d({_al_u1739_o,\t/a/EX_op [4]}),
    .mi({open_n4494,\t/a/EX_op [4]}),
    .sr(rst_pad),
    .f({_al_u1740_o,\t/a/EX_operation [1]}),
    .q({open_n4498,\t/a/MEM_op [4]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*D)"),
    //.LUT1("(~C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110000000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1741|t/a/ex_mem/reg2_b6  (
    .b({\t/a/EX_op [5],\t/a/EX_op [5]}),
    .c({\t/a/EX_op [6],\t/a/EX_op [6]}),
    .clk(clock_pad),
    .d({_al_u1740_o,_al_u1740_o}),
    .mi({open_n4512,\t/a/EX_op [6]}),
    .sr(rst_pad),
    .f({\t/a/aluin/n11_lutinv ,\t/a/aluin/n12_lutinv }),
    .q({open_n4516,\t/a/MEM_op [6]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1744|_al_u1729  (
    .a({\t/a/EX_rd [1],\t/a/MEM_rd [0]}),
    .b({\t/a/EX_rd [3],\t/a/MEM_rd [3]}),
    .c(\t/a/ID_rs1 [1:0]),
    .d({\t/a/ID_rs1 [3],\t/a/ID_rs1 [3]}),
    .f({_al_u1744_o,_al_u1729_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(D*~B)*~(~C*A))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1100010011110101),
    .MODE("LOGIC"))
    \_al_u1745|_al_u1736  (
    .a({\t/a/EX_rd [2],open_n4541}),
    .b({\t/a/EX_rd [3],open_n4542}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs2 [1]}),
    .d({\t/a/ID_rs1 [3],\t/a/EX_rd [1]}),
    .f({_al_u1745_o,_al_u1736_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1746|_al_u1743  (
    .a({_al_u1743_o,_al_u1742_o}),
    .b({_al_u1744_o,\t/a/EX_rd [0]}),
    .c({_al_u1745_o,\t/a/EX_rd [1]}),
    .d({\t/a/EX_rd [4],\t/a/ID_rs1 [0]}),
    .e({\t/a/ID_rs1 [4],\t/a/ID_rs1 [1]}),
    .f({\t/a/risk_jump/n11_lutinv ,_al_u1743_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(0*~(~A*~((~D*~B))*~(C)+~A*(~D*~B)*~(C)+~(~A)*(~D*~B)*C+~A*(~D*~B)*C))"),
    //.LUT1("(1*~(~A*~((~D*~B))*~(C)+~A*(~D*~B)*~(C)+~(~A)*(~D*~B)*C+~A*(~D*~B)*C))"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1111101011001010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1749 (
    .a({_al_u1733_o,_al_u1733_o}),
    .b({\t/a/risk_jump/n35_lutinv ,\t/a/risk_jump/n35_lutinv }),
    .c({\t/a/aluin/n11_lutinv ,\t/a/aluin/n11_lutinv }),
    .d({\t/a/risk_jump/n11_lutinv ,\t/a/risk_jump/n11_lutinv }),
    .mi({open_n4597,\t/a/condition/n1_lutinv }),
    .fx({open_n4602,\t/a/condition/n0_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*~(D*A)))"),
    //.LUT1("(~B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0011001000110000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"))
    \_al_u1758|_al_u1779  (
    .a({\t/a/condition/n5 [31],\t/a/condition/n5 [12]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [31],\t/a/ID_jump_addr [12]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*~(D*A)))"),
    //.LUTF1("(~B*~(~C*~(D*A)))"),
    //.LUTG0("(~B*~(~C*~(D*A)))"),
    //.LUTG1("(~B*~(~C*~(D*A)))"),
    .INIT_LUTF0(16'b0011001000110000),
    .INIT_LUTF1(16'b0011001000110000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0011001000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1759|_al_u1778  (
    .a({\t/a/condition/n5 [30],\t/a/condition/n5 [13]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [30],\t/a/ID_jump_addr [13]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*~(D*A)))"),
    //.LUTF1("(~B*~(~C*~(D*A)))"),
    //.LUTG0("(~B*~(~C*~(D*A)))"),
    //.LUTG1("(~B*~(~C*~(D*A)))"),
    .INIT_LUTF0(16'b0011001000110000),
    .INIT_LUTF1(16'b0011001000110000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0011001000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1761|_al_u1777  (
    .a({\t/a/condition/n5 [29],\t/a/condition/n5 [14]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [29],\t/a/ID_jump_addr [14]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*~(D*A)))"),
    //.LUT1("(~B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0011001000110000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"))
    \_al_u1762|_al_u1776  (
    .a({\t/a/condition/n5 [28],\t/a/condition/n5 [15]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [28],\t/a/ID_jump_addr [15]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*~(D*A)))"),
    //.LUT1("(~B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0011001000110000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"))
    \_al_u1763|_al_u1775  (
    .a({\t/a/condition/n5 [27],\t/a/condition/n5 [16]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [27],\t/a/ID_jump_addr [16]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*~(D*A)))"),
    //.LUTF1("(~B*~(~C*~(D*A)))"),
    //.LUTG0("(~B*~(~C*~(D*A)))"),
    //.LUTG1("(~B*~(~C*~(D*A)))"),
    .INIT_LUTF0(16'b0011001000110000),
    .INIT_LUTF1(16'b0011001000110000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0011001000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1764|_al_u1774  (
    .a({\t/a/condition/n5 [26],\t/a/condition/n5 [17]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [26],\t/a/ID_jump_addr [17]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*~(D*A)))"),
    //.LUTF1("(~B*~(~C*~(D*A)))"),
    //.LUTG0("(~B*~(~C*~(D*A)))"),
    //.LUTG1("(~B*~(~C*~(D*A)))"),
    .INIT_LUTF0(16'b0011001000110000),
    .INIT_LUTF1(16'b0011001000110000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0011001000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1765|_al_u1773  (
    .a({\t/a/condition/n5 [25],\t/a/condition/n5 [18]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [25],\t/a/ID_jump_addr [18]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*~(D*A)))"),
    //.LUT1("(~B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0011001000110000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"))
    \_al_u1766|_al_u1772  (
    .a({\t/a/condition/n5 [24],\t/a/condition/n5 [19]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [24],\t/a/ID_jump_addr [19]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*~(D*A)))"),
    //.LUT1("(~B*~(~C*~(D*A)))"),
    .INIT_LUT0(16'b0011001000110000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"))
    \_al_u1767|_al_u1770  (
    .a({\t/a/condition/n5 [23],\t/a/condition/n5 [20]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f({\t/a/ID_jump_addr [23],\t/a/ID_jump_addr [20]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*~(D*A)))"),
    //.LUTF1("(~B*~(~C*~(D*A)))"),
    //.LUTG0("(~B*~(~C*~(D*A)))"),
    //.LUTG1("(~B*~(~C*~(D*A)))"),
    .INIT_LUTF0(16'b0011001000110000),
    .INIT_LUTF1(16'b0011001000110000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0011001000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1768|_al_u1769  (
    .a(\t/a/condition/n5 [22:21]),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/sel0_b12/B1 ,\t/a/condition/sel0_b12/B1 }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .f(\t/a/ID_jump_addr [22:21]));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUT1("(~B*~(~(1*C)*~(D*A)))"),
    .INIT_LUT0(16'b0010001000000000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1771 (
    .a({\t/a/condition/n5 [2],\t/a/condition/n5 [2]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/n1_lutinv ,\t/a/condition/n1_lutinv }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .mi({open_n4837,\t/a/ID_rd [2]}),
    .fx({open_n4842,\t/a/ID_jump_addr [2]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUT1("(~B*~(~(1*C)*~(D*A)))"),
    .INIT_LUT0(16'b0010001000000000),
    .INIT_LUT1(16'b0011001000110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1780 (
    .a({\t/a/condition/n5 [11],\t/a/condition/n5 [11]}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/n1_lutinv ,\t/a/condition/n1_lutinv }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .mi({open_n4857,\t/a/ID_rd [0]}),
    .fx({open_n4862,\t/a/ID_jump_addr [11]}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1783|t/a/id_ex/reg4_b1  (
    .a({\t/a/MEM_rd [0],\t/a/aluin/sel1_b16/B9 }),
    .b({\t/a/MEM_rd [1],_al_u2007_o}),
    .c({\t/a/EX_rs1 [0],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_rs1 [1],\t/a/EX_rs1 [1]}),
    .mi({open_n4876,\t/a/ID_rs1 [1]}),
    .sr(rst_pad),
    .f({_al_u1783_o,\t/a/EX_B [16]}),
    .q({open_n4880,\t/a/EX_rs1 [1]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~A*~(D*C))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("~(~B*~A*~(D*C))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111011101110),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1111111011101110),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1784|t/a/id_ex/reg4_b4  (
    .a({_al_u1783_o,\t/a/aluin/sel1_b19/B9 }),
    .b({\t/a/MEM_rd [2],_al_u2007_o}),
    .c({\t/a/MEM_rd [4],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_rs1 [2],\t/a/EX_rs1 [4]}),
    .e({\t/a/EX_rs1 [4],open_n4882}),
    .mi({open_n4884,\t/a/ID_rs1 [4]}),
    .sr(rst_pad),
    .f({_al_u1784_o,\t/a/EX_B [19]}),
    .q({open_n4899,\t/a/EX_rs1 [4]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1785|_al_u1727  (
    .c({\t/a/EX_rs1 [1],\t/a/ID_rs1 [1]}),
    .d({\t/a/MEM_rd [1],\t/a/MEM_rd [1]}),
    .f({_al_u1785_o,_al_u1727_o}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~A*~(D*C))"),
    //.LUTF1("(~A*~(0@C)*~(D*~B))"),
    //.LUTG0("~(~B*~A*~(D*C))"),
    //.LUTG1("(~A*~(1@C)*~(D*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111011101110),
    .INIT_LUTF1(16'b0000010000000101),
    .INIT_LUTG0(16'b1111111011101110),
    .INIT_LUTG1(16'b0100000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1786|t/a/id_ex/reg4_b3  (
    .a({_al_u1785_o,\t/a/aluin/sel1_b18/B9 }),
    .b({\t/a/MEM_rd [0],_al_u2007_o}),
    .c({\t/a/MEM_rd [3],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_rs1 [0],\t/a/EX_rs1 [3]}),
    .e({\t/a/EX_rs1 [3],open_n4929}),
    .mi({open_n4931,\t/a/ID_rs1 [3]}),
    .sr(rst_pad),
    .f({_al_u1786_o,\t/a/EX_B [18]}),
    .q({open_n4946,\t/a/EX_rs1 [3]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1787|_al_u1724  (
    .c({_al_u1786_o,\t/a/ID_rs2 [2]}),
    .d({_al_u1784_o,\t/a/MEM_rd [2]}),
    .f({\t/a/n9_lutinv ,_al_u1724_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"))
    \_al_u1788|_al_u328  (
    .a({\t/a/EX_rs1 [3],open_n4975}),
    .b({\t/a/EX_rs1 [4],open_n4976}),
    .c({\t/a/WB_rd [3],\t/a/WB_rd [1]}),
    .d({\t/a/WB_rd [4],\t/a/ID_rs1 [1]}),
    .f({_al_u1788_o,_al_u328_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(0*~C)*~(~D*B))"),
    //.LUT1("(A*~(1*~C)*~(~D*B))"),
    .INIT_LUT0(16'b1010101000100010),
    .INIT_LUT1(16'b1010000000100000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1789 (
    .a({_al_u1788_o,_al_u1788_o}),
    .b({\t/a/EX_rs1 [0],\t/a/EX_rs1 [0]}),
    .c({\t/a/EX_rs1 [1],\t/a/EX_rs1 [1]}),
    .d({\t/a/WB_rd [0],\t/a/WB_rd [0]}),
    .mi({open_n5009,\t/a/WB_rd [1]}),
    .fx({open_n5014,_al_u1789_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"))
    \_al_u1791|_al_u1043  (
    .a({\t/a/EX_rs1 [1],open_n5017}),
    .b({\t/a/EX_rs1 [4],open_n5018}),
    .c({\t/a/WB_rd [1],\t/a/WB_rd [1]}),
    .d({\t/a/WB_rd [4],\t/a/ID_rs2 [1]}),
    .f({_al_u1791_o,_al_u1043_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(C*B*~A*~(0@D))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(C*B*~A*~(1@D))"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b0000000001000000),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b0100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1792|_al_u1790  (
    .a({\t/a/n9_lutinv ,_al_u1789_o}),
    .b({_al_u1790_o,\t/a/EX_rs1 [0]}),
    .c({_al_u1791_o,\t/a/EX_rs1 [3]}),
    .d({\t/a/EX_rs1 [2],\t/a/WB_rd [0]}),
    .e({\t/a/WB_rd [2],\t/a/WB_rd [3]}),
    .f({_al_u1792_o,_al_u1790_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~A*~(D*C*B))"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0001010101010101),
    .MODE("LOGIC"))
    \_al_u1794|_al_u1795  (
    .a({\t/a/regfile/n46 [0],open_n5061}),
    .b({_al_u1793_o,open_n5062}),
    .c({\t/a/WB_op [0],\t/a/n19 }),
    .d({\t/a/WB_op [1],_al_u1792_o}),
    .f({\t/a/n19 ,\t/a/alu_A_select [1]}));
  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*~A)"),
    //.LUTF1("(~A*~(D*C*B))"),
    //.LUTG0("(~1*~D*~C*~B*~A)"),
    //.LUTG1("(~A*~(D*C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0001010101010101),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0001010101010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1797|t/a/mem_wb/reg2_b4  (
    .a({_al_u1796_o,\t/a/MEM_rd [0]}),
    .b({_al_u251_o,\t/a/MEM_rd [1]}),
    .c({_al_u252_o,\t/a/MEM_rd [2]}),
    .clk(clock_pad),
    .d({\t/a/MEM_op [5],\t/a/MEM_rd [3]}),
    .e({open_n5084,\t/a/MEM_rd [4]}),
    .mi({open_n5086,\t/a/MEM_rd [4]}),
    .sr(rst_pad),
    .f({_al_u1797_o,_al_u1796_o}),
    .q({open_n5101,\t/a/WB_rd [4]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~B*~D))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*~(~B*~D))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111000011000000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111000011000000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1798|_al_u1733  (
    .b({open_n5104,\t/a/risk_jump/n24_lutinv }),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .d({_al_u1797_o,\t/a/risk_jump/n42_lutinv }),
    .f({_al_u1798_o,_al_u1733_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1800|t/a/regfile/reg0_b105  (
    .a({\t/a/alu_A_select [1],_al_u2606_o}),
    .b({\t/a/alu_A_select [0],_al_u2610_o}),
    .c({\t/a/MEM_aludat [9],\t/a/MEM_aludat [9]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [9],\t/a/reg_writedat [9]}),
    .mi({open_n5139,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u1800_o,_al_u2716_o}),
    .q({open_n5143,\t/a/regfile/regfile$3$ [9]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(~C*B))"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("(~D*~(~C*B))"),
    //.LUTG1("(D*C*~B*A)"),
    .INIT_LUTF0(16'b0000000011110011),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b0000000011110011),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1802|_al_u1806  (
    .a({_al_u1801_o,open_n5144}),
    .b({\t/a/EX_op [4],_al_u1803_o}),
    .c({\t/a/EX_op [5],\t/a/EX_op [5]}),
    .d({\t/a/EX_op [6],_al_u1802_o}),
    .f({_al_u1802_o,_al_u1806_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u1804|_al_u1114  (
    .a({open_n5169,\t/a/ID_rs2 [0]}),
    .b({open_n5170,\t/a/ID_rs2 [1]}),
    .c({_al_u1803_o,\t/a/regfile/regfile$6$ [6]}),
    .d({_al_u1802_o,\t/a/regfile/regfile$7$ [6]}),
    .f({\t/a/aluin/n5_lutinv ,_al_u1114_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1807|t/a/regfile/reg0_b169  (
    .a({open_n5191,_al_u1800_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [9],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b9/B0 ,\t/a/reg_writedat [9]}),
    .mi({open_n5202,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [9],\t/a/aluin/sel0_b9/B0 }),
    .q({open_n5206,\t/a/regfile/regfile$5$ [9]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1808|t/a/regfile/reg0_b104  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [8],\t/a/MEM_aludat [8]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [8],\t/a/reg_writedat [8]}),
    .mi({open_n5217,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u1808_o,_al_u2722_o}),
    .q({open_n5221,\t/a/regfile/regfile$3$ [8]}));  // register.v(63)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTG1("~(~D*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111100010),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b1111001111100010),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1810|t/a/id_ex/reg7_b8  (
    .a({open_n5222,_al_u2807_o}),
    .b({_al_u1806_o,\t/a/condition/n0_lutinv }),
    .c({\t/a/EX_memstraddr [8],\t/a/ID_memstraddr [8]}),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b8/B0 ,\t/memstraddress [8]}),
    .mi({open_n5227,\t/a/ID_memstraddr [8]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [8],_al_u2815_o}),
    .q({open_n5242,\t/a/EX_memstraddr [8]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG0("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT_LUTF0(16'b0000010000010101),
    .INIT_LUTF1(16'b0000010000010101),
    .INIT_LUTG0(16'b0000010000010101),
    .INIT_LUTG1(16'b0000010000010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1811|_al_u1817  (
    .a({\t/a/alu_A_select [1],\t/a/alu_A_select [1]}),
    .b({\t/a/alu_A_select [0],\t/a/alu_A_select [0]}),
    .c({\t/a/MEM_aludat [7],\t/a/MEM_aludat [5]}),
    .d({\t/a/EX_regdat1 [7],\t/a/EX_regdat1 [5]}),
    .f({_al_u1811_o,_al_u1817_o}));
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1814|t/a/if_id/reg5_b6  (
    .a({\t/a/alu_A_select [1],open_n5267}),
    .b({\t/a/alu_A_select [0],\t/a/MEM_aludat [6]}),
    .c({\t/a/MEM_aludat [6],\t/memstraddress [6]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [6],\t/busarbitration/n3 }),
    .mi({open_n5278,\t/memstraddress [6]}),
    .sr(rst_pad),
    .f({_al_u1814_o,addr[6]}),
    .q({open_n5282,\t/a/ID_memstraddr [6]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUT1("~(~D*~(C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111100010),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1819|t/a/id_ex/reg7_b5  (
    .a({open_n5283,_al_u2807_o}),
    .b({_al_u1806_o,\t/a/condition/n0_lutinv }),
    .c({\t/a/EX_memstraddr [5],\t/a/ID_memstraddr [5]}),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b5/B0 ,\t/memstraddress [5]}),
    .mi({open_n5295,\t/a/ID_memstraddr [5]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [5],_al_u2822_o}),
    .q({open_n5299,\t/a/EX_memstraddr [5]}));  // flow_line_reg.v(139)
  EG_PHY_PAD #(
    //.LOCATION("P161"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u182 (
    .ipad(clock),
    .di(clock_pad));  // __top.v(4)
  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~A*~(D*~B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000101),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1820|t/a/ex_mem/reg4_b4  (
    .a({\t/a/alu_A_select [1],_al_u2541_o}),
    .b({\t/a/alu_A_select [0],\t/a/alu/n6 [4]}),
    .c({\t/a/MEM_aludat [4],_al_u2547_o}),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [4],_al_u2126_o}),
    .sr(rst_pad),
    .f({_al_u1820_o,\t/a/aludat [4]}),
    .q({open_n5333,\t/a/MEM_aludat [4]}));  // flow_line_reg.v(191)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1823|t/a/regfile/reg0_b1023  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [31],\t/a/MEM_aludat [31]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [31],\t/a/reg_writedat [31]}),
    .mi({open_n5344,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1823_o,_al_u2617_o}),
    .q({open_n5348,\t/a/regfile/regfile$31$ [31]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1826|t/a/regfile/reg0_b1022  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [30],\t/a/MEM_aludat [30]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [30],\t/a/reg_writedat [30]}),
    .mi({open_n5359,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1826_o,_al_u2621_o}),
    .q({open_n5363,\t/a/regfile/regfile$31$ [30]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1828|t/a/regfile/reg0_b190  (
    .a({open_n5364,_al_u1826_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [30],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b30/B0 ,\t/a/reg_writedat [30]}),
    .mi({open_n5375,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [30],\t/a/aluin/sel0_b30/B0 }),
    .q({open_n5379,\t/a/regfile/regfile$5$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT_LUTF0(16'b0000010010001100),
    .INIT_LUTF1(16'b0000010000010101),
    .INIT_LUTG0(16'b0000010010001100),
    .INIT_LUTG1(16'b0000010000010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1829|_al_u461  (
    .a({\t/a/alu_A_select [1],\t/a/ID_rs1 [0]}),
    .b({\t/a/alu_A_select [0],\t/a/ID_rs1 [1]}),
    .c({\t/a/MEM_aludat [3],\t/a/regfile/regfile$6$ [3]}),
    .d({\t/a/EX_regdat1 [3],\t/a/regfile/regfile$7$ [3]}),
    .f({_al_u1829_o,_al_u461_o}));
  EG_PHY_PAD #(
    //.LOCATION("P136"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u183 (
    .ipad(rst),
    .di(rst_pad));  // __top.v(3)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1832|t/a/regfile/reg0_b1021  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [29],\t/a/MEM_aludat [29]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [29],\t/a/reg_writedat [29]}),
    .mi({open_n5431,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1832_o,_al_u2625_o}),
    .q({open_n5435,\t/a/regfile/regfile$31$ [29]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1834|t/a/regfile/reg0_b189  (
    .a({open_n5436,_al_u1832_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [29],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b29/B0 ,\t/a/reg_writedat [29]}),
    .mi({open_n5447,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [29],\t/a/aluin/sel0_b29/B0 }),
    .q({open_n5451,\t/a/regfile/regfile$5$ [29]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1835|t/a/regfile/reg0_b1020  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [28],\t/a/MEM_aludat [28]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [28],\t/a/reg_writedat [28]}),
    .mi({open_n5462,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1835_o,_al_u2629_o}),
    .q({open_n5466,\t/a/regfile/regfile$31$ [28]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1838|t/a/regfile/reg0_b1019  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [27],\t/a/MEM_aludat [27]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [27],\t/a/reg_writedat [27]}),
    .mi({open_n5477,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1838_o,_al_u2633_o}),
    .q({open_n5481,\t/a/regfile/regfile$31$ [27]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1841|t/a/regfile/reg0_b1018  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [26],\t/a/MEM_aludat [26]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [26],\t/a/reg_writedat [26]}),
    .mi({open_n5492,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1841_o,_al_u2637_o}),
    .q({open_n5496,\t/a/regfile/regfile$31$ [26]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1843|t/a/regfile/reg0_b186  (
    .a({open_n5497,_al_u1841_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [26],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b26/B0 ,\t/a/reg_writedat [26]}),
    .mi({open_n5508,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [26],\t/a/aluin/sel0_b26/B0 }),
    .q({open_n5512,\t/a/regfile/regfile$5$ [26]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1844|t/a/regfile/reg0_b1017  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [25],\t/a/MEM_aludat [25]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [25],\t/a/reg_writedat [25]}),
    .mi({open_n5523,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1844_o,_al_u2641_o}),
    .q({open_n5527,\t/a/regfile/regfile$31$ [25]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1846|t/a/regfile/reg0_b185  (
    .a({open_n5528,_al_u1844_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [25],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b25/B0 ,\t/a/reg_writedat [25]}),
    .mi({open_n5539,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [25],\t/a/aluin/sel0_b25/B0 }),
    .q({open_n5543,\t/a/regfile/regfile$5$ [25]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1847|t/a/regfile/reg0_b1016  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [24],\t/a/MEM_aludat [24]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [24],\t/a/reg_writedat [24]}),
    .mi({open_n5554,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1847_o,_al_u2645_o}),
    .q({open_n5558,\t/a/regfile/regfile$31$ [24]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1849|t/a/regfile/reg0_b184  (
    .a({open_n5559,_al_u1847_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [24],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b24/B0 ,\t/a/reg_writedat [24]}),
    .mi({open_n5563,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [24],\t/a/aluin/sel0_b24/B0 }),
    .q({open_n5578,\t/a/regfile/regfile$5$ [24]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1850|t/a/regfile/reg0_b1015  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [23],\t/a/MEM_aludat [23]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [23],\t/a/reg_writedat [23]}),
    .mi({open_n5589,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1850_o,_al_u2649_o}),
    .q({open_n5593,\t/a/regfile/regfile$31$ [23]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1852|t/a/regfile/reg0_b183  (
    .a({open_n5594,_al_u1850_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [23],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b23/B0 ,\t/a/reg_writedat [23]}),
    .mi({open_n5598,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [23],\t/a/aluin/sel0_b23/B0 }),
    .q({open_n5613,\t/a/regfile/regfile$5$ [23]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1853|t/a/regfile/reg0_b1014  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [22],\t/a/MEM_aludat [22]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [22],\t/a/reg_writedat [22]}),
    .mi({open_n5624,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1853_o,_al_u2653_o}),
    .q({open_n5628,\t/a/regfile/regfile$31$ [22]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1856|t/a/regfile/reg0_b1013  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [21],\t/a/MEM_aludat [21]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [21],\t/a/reg_writedat [21]}),
    .mi({open_n5639,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1856_o,_al_u2657_o}),
    .q({open_n5643,\t/a/regfile/regfile$31$ [21]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1859|t/a/regfile/reg0_b1012  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [20],\t/a/MEM_aludat [20]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [20],\t/a/reg_writedat [20]}),
    .mi({open_n5654,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1859_o,_al_u2661_o}),
    .q({open_n5658,\t/a/regfile/regfile$31$ [20]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1861|t/a/regfile/reg0_b180  (
    .a({open_n5659,_al_u1859_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [20],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b20/B0 ,\t/a/reg_writedat [20]}),
    .mi({open_n5663,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [20],\t/a/aluin/sel0_b20/B0 }),
    .q({open_n5678,\t/a/regfile/regfile$5$ [20]}));  // register.v(63)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1862|t/a/id_ex/reg8_b2  (
    .a({\t/a/alu_A_select [1],_al_u333_o}),
    .b({\t/a/alu_A_select [0],_al_u532_o}),
    .c({\t/a/MEM_aludat [2],_al_u542_o}),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [2],\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u1862_o,\t/a/ID_read_dat1 [2]}),
    .q({open_n5695,\t/a/EX_regdat1 [2]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("~(~D*~(C*~B))"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"))
    \_al_u1864|_al_u1241  (
    .a({open_n5696,\t/a/ID_rs2 [0]}),
    .b({_al_u1806_o,\t/a/ID_rs2 [1]}),
    .c({\t/a/EX_memstraddr [2],\t/a/regfile/regfile$0$ [2]}),
    .d({\t/a/aluin/sel0_b2/B0 ,\t/a/regfile/regfile$1$ [2]}),
    .f({\t/a/EX_A [2],_al_u1241_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1865|t/a/regfile/reg0_b1011  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [19],\t/a/MEM_aludat [19]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [19],\t/a/reg_writedat [19]}),
    .mi({open_n5727,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1865_o,_al_u2665_o}),
    .q({open_n5731,\t/a/regfile/regfile$31$ [19]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1868|t/a/regfile/reg0_b1010  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [18],\t/a/MEM_aludat [18]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [18],\t/a/reg_writedat [18]}),
    .mi({open_n5742,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1868_o,_al_u2669_o}),
    .q({open_n5746,\t/a/regfile/regfile$31$ [18]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1871|t/a/regfile/reg0_b1009  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [17],\t/a/MEM_aludat [17]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [17],\t/a/reg_writedat [17]}),
    .mi({open_n5757,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1871_o,_al_u2673_o}),
    .q({open_n5761,\t/a/regfile/regfile$31$ [17]}));  // register.v(63)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1874|t/a/id_ex/reg8_b16  (
    .a({\t/a/alu_A_select [1],_al_u333_o}),
    .b({\t/a/alu_A_select [0],_al_u847_o}),
    .c({\t/a/MEM_aludat [16],_al_u857_o}),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [16],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1874_o,\t/a/ID_read_dat1 [16]}),
    .q({open_n5778,\t/a/EX_regdat1 [16]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~B))"),
    //.LUT1("~(~D*~(C*~B))"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"))
    \_al_u1876|_al_u1891  (
    .b({_al_u1806_o,_al_u1806_o}),
    .c({\t/a/EX_memstraddr [16],\t/a/EX_memstraddr [11]}),
    .d({\t/a/aluin/sel0_b16/B0 ,\t/a/aluin/sel0_b11/B0 }),
    .f({\t/a/EX_A [16],\t/a/EX_A [11]}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1877|t/a/regfile/reg0_b655  (
    .a({\t/a/alu_A_select [1],\t/a/ID_rs1 [0]}),
    .b({\t/a/alu_A_select [0],\t/a/ID_rs1 [1]}),
    .c({\t/a/MEM_aludat [15],\t/a/regfile/regfile$20$ [15]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [15],\t/a/regfile/regfile$21$ [15]}),
    .mi({open_n5811,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1877_o,_al_u869_o}),
    .q({open_n5815,\t/a/regfile/regfile$20$ [15]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~B*A)"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(~D*C*~B*A)"),
    //.LUTG1("~(~D*~(C*~B))"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1879|_al_u1803  (
    .a({open_n5816,_al_u1801_o}),
    .b({_al_u1806_o,\t/a/EX_op [3]}),
    .c({\t/a/EX_memstraddr [15],\t/a/EX_op [4]}),
    .d({\t/a/aluin/sel0_b15/B0 ,\t/a/EX_op [6]}),
    .f({\t/a/EX_A [15],_al_u1803_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1880|t/a/regfile/reg0_b1006  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [14],\t/a/MEM_aludat [14]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [14],\t/a/reg_writedat [14]}),
    .mi({open_n5851,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1880_o,_al_u2693_o}),
    .q({open_n5855,\t/a/regfile/regfile$31$ [14]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1882|t/a/regfile/reg0_b142  (
    .a({open_n5856,_al_u1880_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [14],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b14/B0 ,\t/a/reg_writedat [14]}),
    .mi({open_n5860,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [14],\t/a/aluin/sel0_b14/B0 }),
    .q({open_n5875,\t/a/regfile/regfile$4$ [14]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1883|t/a/regfile/reg0_b1005  (
    .a({\t/a/alu_A_select [1],_al_u2614_o}),
    .b({\t/a/alu_A_select [0],_al_u2616_o}),
    .c({\t/a/MEM_aludat [13],\t/a/MEM_aludat [13]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [13],\t/a/reg_writedat [13]}),
    .mi({open_n5886,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1883_o,_al_u2697_o}),
    .q({open_n5890,\t/a/regfile/regfile$31$ [13]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1885|t/a/regfile/reg0_b141  (
    .a({open_n5891,_al_u1883_o}),
    .b({_al_u1806_o,\t/a/alu_A_select [1]}),
    .c({\t/a/EX_memstraddr [13],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel0_b13/B0 ,\t/a/reg_writedat [13]}),
    .mi({open_n5895,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({\t/a/EX_A [13],\t/a/aluin/sel0_b13/B0 }),
    .q({open_n5910,\t/a/regfile/regfile$4$ [13]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1886|t/a/regfile/reg0_b140  (
    .a({\t/a/alu_A_select [1],_al_u1886_o}),
    .b({\t/a/alu_A_select [0],\t/a/alu_A_select [1]}),
    .c({\t/a/MEM_aludat [12],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [12],\t/a/reg_writedat [12]}),
    .mi({open_n5921,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1886_o,\t/a/aluin/sel0_b12/B0 }),
    .q({open_n5925,\t/a/regfile/regfile$4$ [12]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1889|t/a/regfile/reg0_b139  (
    .a({\t/a/alu_A_select [1],_al_u1889_o}),
    .b({\t/a/alu_A_select [0],\t/a/alu_A_select [1]}),
    .c({\t/a/MEM_aludat [11],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [11],\t/a/reg_writedat [11]}),
    .mi({open_n5936,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u1889_o,\t/a/aluin/sel0_b11/B0 }),
    .q({open_n5940,\t/a/regfile/regfile$4$ [11]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b0000010000010101),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000010000010101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1892|t/a/regfile/reg0_b138  (
    .a({\t/a/alu_A_select [1],_al_u1892_o}),
    .b({\t/a/alu_A_select [0],\t/a/alu_A_select [1]}),
    .c({\t/a/MEM_aludat [10],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [10],\t/a/reg_writedat [10]}),
    .mi({open_n5944,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1892_o,\t/a/aluin/sel0_b10/B0 }),
    .q({open_n5959,\t/a/regfile/regfile$4$ [10]}));  // register.v(63)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1895|t/a/id_ex/reg8_b1  (
    .a({\t/a/alu_A_select [1],_al_u333_o}),
    .b({\t/a/alu_A_select [0],_al_u763_o}),
    .c({\t/a/MEM_aludat [1],_al_u773_o}),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [1],\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u1895_o,\t/a/ID_read_dat1 [1]}),
    .q({open_n5976,\t/a/EX_regdat1 [1]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("~(~D*~(C*~B))"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"))
    \_al_u1897|_al_u2217  (
    .b({_al_u1806_o,open_n5979}),
    .c({\t/a/EX_memstraddr [1],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel0_b1/B0 ,\t/a/alu/n170_lutinv }),
    .f({\t/a/EX_A [1],\t/a/alu/n202_lutinv }));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010000010101),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1898|t/a/regfile/reg0_b992  (
    .a({\t/a/alu_A_select [1],_al_u2606_o}),
    .b({\t/a/alu_A_select [0],_al_u2610_o}),
    .c({\t/a/MEM_aludat [0],\t/a/MEM_aludat [0]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_regdat1 [0],\t/a/reg_writedat [0]}),
    .mi({open_n6010,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u1898_o,_al_u2758_o}),
    .q({open_n6014,\t/a/regfile/regfile$31$ [0]}));  // register.v(63)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~B))"),
    //.LUTF1("(C*~A*~(~D*B))"),
    //.LUTG0("~(~D*~(C*~B))"),
    //.LUTG1("(C*~A*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100110000),
    .INIT_LUTF1(16'b0101000000010000),
    .INIT_LUTG0(16'b1111111100110000),
    .INIT_LUTG1(16'b0101000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1899|t/a/id_ex/reg7_b0  (
    .a({_al_u1898_o,open_n6015}),
    .b({\t/a/alu_A_select [1],_al_u1806_o}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/EX_memstraddr [0]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [0],\t/a/aluin/sel0_b0/B0 }),
    .mi({open_n6020,\t/a/ID_memstraddr [0]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b0/B0 ,\t/a/EX_A [0]}),
    .q({open_n6035,\t/a/EX_memstraddr [0]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUTG1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111001001010000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0111001001010000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1901|t/a/mem_wb/reg0_b7  (
    .a({open_n6036,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({open_n6037,_al_u1908_o}),
    .c({i_data[7],\t/a/MEM_aludat [7]}),
    .clk(clock_pad),
    .d({\t/busarbitration/mux5_b0_sel_is_3_o ,i_data[7]}),
    .sr(rst_pad),
    .f({\t/a/mux4_b7/B0_0 ,open_n6055}),
    .q({open_n6059,\t/a/reg_writedat [7]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*B*A*(D@C))"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("(~1*B*A*(D@C))"),
    //.LUTG1("(~D*~C*~B*A)"),
    .INIT_LUTF0(16'b0000100010000000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1902|_al_u1027  (
    .a({\t/a/mux4_b7/B0_0 ,memwrite_cs}),
    .b({\t/a/MEM_fun3 [0],\t/a/MEM_regdat2 [13]}),
    .c(\t/a/MEM_fun3 [1:0]),
    .d(\t/a/MEM_fun3 [2:1]),
    .e({open_n6062,\t/a/MEM_fun3 [2]}),
    .f({_al_u1902_o,o_data[13]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*C*~B*A)"),
    //.LUTF1("(~(D)*~(B)*~(C)+D*B*~(C)+~(D)*~(B)*C+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~D*C*~B*A)"),
    //.LUTG1("(~(D)*~(B)*~(C)+D*B*~(C)+~(D)*~(B)*C+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b1100110011110011),
    .INIT_LUTG0(16'b0000000000100000),
    .INIT_LUTG1(16'b1100110011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1903|_al_u1918  (
    .a({open_n6083,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b(\t/a/MEM_fun3 [1:0]),
    .c(\t/a/MEM_fun3 [2:1]),
    .d({\t/a/MEM_fun3 [0],\t/a/MEM_fun3 [2]}),
    .f({_al_u1903_o,_al_u1918_o}));
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1904|t/a/if_id/reg2_b2  (
    .a({open_n6108,\t/a/if_id/n9 }),
    .b({_al_u1903_o,\t/busarbitration/n3 }),
    .c({i_data[9],\t/busarbitration/instruction [9]}),
    .clk(clock_pad),
    .d({\t/busarbitration/mux5_b0_sel_is_3_o ,i_data[9]}),
    .sr(rst_pad),
    .f({_al_u1904_o,open_n6126}),
    .q({open_n6130,\t/a/ID_rd [2]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1906|t/a/if_id/reg2_b1  (
    .a({open_n6131,\t/a/if_id/n9 }),
    .b({_al_u1903_o,\t/busarbitration/n3 }),
    .c({i_data[8],\t/busarbitration/instruction [8]}),
    .clk(clock_pad),
    .d({\t/busarbitration/mux5_b0_sel_is_3_o ,i_data[8]}),
    .sr(rst_pad),
    .f({_al_u1906_o,open_n6149}),
    .q({open_n6153,\t/a/ID_rd [1]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*B*D)"),
    //.LUTF1("(B*~(~C*~D))"),
    //.LUTG0("(~C*B*D)"),
    //.LUTG1("(B*~(~C*~D))"),
    .INIT_LUTF0(16'b0000110000000000),
    .INIT_LUTF1(16'b1100110011000000),
    .INIT_LUTG0(16'b0000110000000000),
    .INIT_LUTG1(16'b1100110011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1908|_al_u1917  (
    .b({\t/a/MEM_fun3 [1],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .c({\t/a/MEM_fun3 [2],\t/a/MEM_fun3 [2]}),
    .d({\t/a/MEM_fun3 [0],_al_u1916_o}),
    .f({_al_u1908_o,_al_u1917_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*A*(~(B)*C*~(D)+B*~(C)*D))"),
    //.LUTF1("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(1*A*(~(B)*C*~(D)+B*~(C)*D))"),
    //.LUTG1("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0011001000010000),
    .INIT_LUTG0(16'b0000100000100000),
    .INIT_LUTG1(16'b0011001000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1916|_al_u1935  (
    .a({\t/a/MEM_fun3 [0],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b(\t/a/MEM_fun3 [1:0]),
    .c({i_data[7],\t/a/MEM_fun3 [1]}),
    .d({i_data[15],\t/a/MEM_fun3 [2]}),
    .e({open_n6182,i_data[15]}),
    .f({_al_u1916_o,_al_u1935_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(~C*~B))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000011111100),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u1940|_al_u2596  (
    .b({open_n6205,i_data[10]}),
    .c({i_data[11],i_data[12]}),
    .d({_al_u1903_o,_al_u1903_o}),
    .f({_al_u1940_o,_al_u2596_o}));
  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111001001010000),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0111001001010000),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1945|t/a/mem_wb/reg0_b3  (
    .a({open_n6226,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({\t/busarbitration/instruction [3],_al_u1908_o}),
    .c({i_data[3],\t/a/MEM_aludat [3]}),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,i_data[3]}),
    .sr(rst_pad),
    .f({\t/instruction$3$_neg_lutinv ,open_n6244}),
    .q({open_n6248,\t/a/reg_writedat [3]}));  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111001001010000),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1946|t/a/mem_wb/reg0_b4  (
    .a({open_n6249,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({\t/busarbitration/instruction [4],_al_u1908_o}),
    .c({i_data[4],\t/a/MEM_aludat [4]}),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,i_data[4]}),
    .sr(rst_pad),
    .f({\t/instruction$4$_neg_lutinv ,open_n6263}),
    .q({open_n6267,\t/a/reg_writedat [4]}));  // flow_line_reg.v(234)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1947|t/a/if_id/reg6_b4  (
    .b({\t/instruction$3$_neg_lutinv ,open_n6270}),
    .c({\t/instruction$4$_neg_lutinv ,\t/instruction$4$_neg_lutinv }),
    .clk(clock_pad),
    .d({_al_u1944_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({_al_u1947_o,open_n6284}),
    .q({open_n6288,\t/a/ID_op [4]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("~((C*B)*~((0*D))*~(A)+(C*B)*(0*D)*~(A)+~((C*B))*(0*D)*A+(C*B)*(0*D)*A)"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("~((C*B)*~((1*D))*~(A)+(C*B)*(1*D)*~(A)+~((C*B))*(1*D)*A+(C*B)*(1*D)*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b1011111110111111),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010110111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1948|t/a/if_id/reg6_b1  (
    .a({\t/busarbitration/n3 ,\t/a/if_id/n9 }),
    .b({\t/busarbitration/instruction [0],\t/busarbitration/n3 }),
    .c({\t/busarbitration/instruction [1],\t/busarbitration/instruction [1]}),
    .clk(clock_pad),
    .d({i_data[1],i_data[1]}),
    .e({i_data[0],open_n6290}),
    .sr(rst_pad),
    .f({_al_u1948_o,open_n6305}),
    .q({open_n6309,\t/a/ID_op [1]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111001001010000),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0111001001010000),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1949|t/a/mem_wb/reg0_b2  (
    .a({open_n6310,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({\t/busarbitration/instruction [2],_al_u1908_o}),
    .c({i_data[2],\t/a/MEM_aludat [2]}),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,i_data[2]}),
    .sr(rst_pad),
    .f({\t/instruction$2$_neg_lutinv ,open_n6328}),
    .q({open_n6332,\t/a/reg_writedat [2]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*~(D*~C*~B*A))"),
    //.LUTF1("(~C*~B*D)"),
    //.LUTG0("(1*~(D*~C*~B*A))"),
    //.LUTG1("(~C*~B*D)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000001100000000),
    .INIT_LUTG0(16'b1111110111111111),
    .INIT_LUTG1(16'b0000001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1950|_al_u2805  (
    .a({open_n6333,_al_u2802_o}),
    .b({_al_u1948_o,_al_u1948_o}),
    .c({\t/instruction$2$_neg_lutinv ,_al_u1944_o}),
    .d({_al_u1947_o,\t/instruction$4$_neg_lutinv }),
    .e({open_n6336,\t/a/n0_lutinv }),
    .f({_al_u1950_o,\t/a/n2 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1010100000100000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1951|_al_u1955  (
    .a({_al_u1950_o,_al_u1950_o}),
    .b({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .c({\t/busarbitration/instruction [29],\t/busarbitration/instruction [25]}),
    .d({i_data[29],i_data[25]}),
    .f({\t/a/IF_skip_addr [9],\t/a/IF_skip_addr [5]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(B*(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUTF0(16'b1010111010101010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1110111011101010),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1952|_al_u2083  (
    .a({_al_u1950_o,_al_u2078_o}),
    .b({\t/busarbitration/n3 ,_al_u2080_o}),
    .c({\t/busarbitration/instruction [28],\t/busarbitration/n3 }),
    .d({i_data[28],\t/busarbitration/instruction [28]}),
    .e({open_n6383,i_data[28]}),
    .f({\t/a/IF_skip_addr [8],\t/a/IF_skip_addr [28]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("~(~A*~(B*(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT_LUTF0(16'b1010111010101010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1110111011101010),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1953|_al_u2084  (
    .a({_al_u1950_o,_al_u2078_o}),
    .b({\t/busarbitration/n3 ,_al_u2080_o}),
    .c({\t/busarbitration/instruction [27],\t/busarbitration/n3 }),
    .d({i_data[27],\t/busarbitration/instruction [27]}),
    .e({open_n6406,i_data[27]}),
    .f({\t/a/IF_skip_addr [7],\t/a/IF_skip_addr [27]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~C*B*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(~C*B*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b1111001111111111),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b1111001111111111),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1956|_al_u289  (
    .b({\t/busarbitration/instruction [24],_al_u252_o}),
    .c({i_data[24],\t/a/MEM_op [6]}),
    .d({\t/busarbitration/n3 ,_al_u251_o}),
    .f({_al_u1956_o,\t/busarbitration/n3 }));
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1957|t/a/if_id/reg4_b4  (
    .c({_al_u1956_o,_al_u1956_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [4],open_n6474}),
    .q({open_n6478,\t/a/ID_rs2 [4]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1959|t/a/if_id/reg4_b3  (
    .c({_al_u1958_o,_al_u1958_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [3],open_n6496}),
    .q({open_n6500,\t/a/ID_rs2 [3]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1960|_al_u2117  (
    .b({\t/busarbitration/instruction [22],\t/busarbitration/instruction [16]}),
    .c({i_data[22],i_data[16]}),
    .d({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .f({_al_u1960_o,_al_u2117_o}));
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1961|t/a/if_id/reg4_b2  (
    .c({_al_u1960_o,_al_u1960_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [2],open_n6544}),
    .q({open_n6548,\t/a/ID_rs2 [2]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1963|t/a/if_id/reg4_b0  (
    .c({_al_u1962_o,_al_u1962_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [11],open_n6566}),
    .q({open_n6570,\t/a/ID_rs2 [0]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1966|t/a/if_id/reg4_b1  (
    .c({_al_u1965_o,_al_u1965_o}),
    .clk(clock_pad),
    .d({_al_u1950_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [1],open_n6588}),
    .q({open_n6592,\t/a/ID_rs2 [1]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1967|t/a/id_ex/reg3_b3  (
    .a({open_n6593,\t/a/aluin/sel1_b23/B9 }),
    .b({open_n6594,_al_u2007_o}),
    .c({\t/a/EX_rs2 [3],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_rd [3],\t/a/EX_rs2 [3]}),
    .mi({open_n6606,\t/a/ID_rs2 [3]}),
    .sr(rst_pad),
    .f({_al_u1967_o,\t/a/EX_B [23]}),
    .q({open_n6610,\t/a/EX_rs2 [3]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u1972|_al_u1978  (
    .c({\t/a/n24_lutinv ,\t/a/n24_lutinv }),
    .d({_al_u1798_o,\t/a/n29 }),
    .f({\t/a/alu_B_select [0],\t/a/alu_B_select [1]}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1973|t/a/id_ex/reg3_b0  (
    .a({open_n6635,\t/a/aluin/n12_lutinv }),
    .b({open_n6636,_al_u1984_o}),
    .c({\t/a/WB_rd [0],\t/a/EX_rs2 [0]}),
    .clk(clock_pad),
    .d({\t/a/EX_rs2 [0],\t/a/EX_rd [0]}),
    .mi({open_n6648,\t/a/ID_rs2 [0]}),
    .sr(rst_pad),
    .f({_al_u1973_o,_al_u2076_o}),
    .q({open_n6652,\t/a/EX_rs2 [0]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0@C)*~(D*~B))"),
    //.LUT1("(~A*~(1@C)*~(D*~B))"),
    .INIT_LUT0(16'b0000010000000101),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1974 (
    .a({_al_u1973_o,_al_u1973_o}),
    .b({\t/a/EX_rs2 [1],\t/a/EX_rs2 [1]}),
    .c({\t/a/EX_rs2 [3],\t/a/EX_rs2 [3]}),
    .d({\t/a/WB_rd [1],\t/a/WB_rd [1]}),
    .mi({open_n6665,\t/a/WB_rd [3]}),
    .fx({open_n6670,_al_u1974_o}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1975|t/a/id_ex/reg3_b1  (
    .a({open_n6673,\t/a/aluin/sel1_b21/B9 }),
    .b({open_n6674,_al_u2007_o}),
    .c({\t/a/WB_rd [1],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_rs2 [1],\t/a/EX_rs2 [1]}),
    .mi({open_n6686,\t/a/ID_rs2 [1]}),
    .sr(rst_pad),
    .f({_al_u1975_o,\t/a/EX_B [21]}),
    .q({open_n6690,\t/a/EX_rs2 [1]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1977|_al_u1976  (
    .a({\t/a/n19 ,_al_u1975_o}),
    .b({_al_u1974_o,\t/a/EX_rs2 [0]}),
    .c({_al_u1976_o,\t/a/EX_rs2 [4]}),
    .d({\t/a/EX_rs2 [2],\t/a/WB_rd [0]}),
    .e({\t/a/WB_rd [2],\t/a/WB_rd [4]}),
    .f({\t/a/n29 ,_al_u1976_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1983|_al_u491  (
    .a({open_n6713,\t/a/ID_rs1 [0]}),
    .b({open_n6714,\t/a/ID_rs1 [1]}),
    .c({\t/a/aluin/n12_lutinv ,\t/a/regfile/regfile$4$ [31]}),
    .d({\t/a/aluin/n11_lutinv ,\t/a/regfile/regfile$5$ [31]}),
    .f({_al_u1983_o,_al_u491_o}));
  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~B*~(D*A)))"),
    //.LUTF1("(A*~(B*~(~D*C)))"),
    //.LUTG0("(C*~(~B*~(D*A)))"),
    //.LUTG1("(A*~(B*~(~D*C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1110000011000000),
    .INIT_LUTF1(16'b0010001010100010),
    .INIT_LUTG0(16'b1110000011000000),
    .INIT_LUTG1(16'b0010001010100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1985|t/a/ex_mem/reg3_b0  (
    .a({_al_u1983_o,_al_u1984_o}),
    .b({_al_u1984_o,\t/a/aluin/n10_lutinv }),
    .c({\t/a/EX_fun3 [0],\t/a/EX_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/EX_fun3 [1],\t/a/EX_op [4]}),
    .mi({open_n6743,\t/a/EX_fun3 [0]}),
    .sr(rst_pad),
    .f({_al_u1985_o,\t/a/EX_operation [0]}),
    .q({open_n6758,\t/a/MEM_fun3 [0]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~D*(B@A)))"),
    //.LUT1("~(~D*~(C*~B))"),
    .INIT_LUT0(16'b1111000010010000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"))
    \_al_u1986|_al_u2495  (
    .a({open_n6759,\t/a/EX_A [9]}),
    .b({_al_u1985_o,\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_fun7 [4],_al_u2431_o}),
    .d({\t/a/aluin/sel1_b9/B9 ,\t/a/EX_operation [0]}),
    .f({\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ,_al_u2495_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1989|t/a/regfile/reg0_b168  (
    .a({open_n6780,_al_u1987_o}),
    .b({_al_u1985_o,\t/a/alu_B_select [1]}),
    .c({\t/a/EX_fun7 [3],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b8/B9 ,\t/a/reg_writedat [8]}),
    .mi({open_n6784,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b8/B9 }),
    .q({open_n6799,\t/a/regfile/regfile$5$ [8]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1992|t/a/regfile/reg0_b167  (
    .a({open_n6800,_al_u1990_o}),
    .b({_al_u1985_o,\t/a/alu_B_select [1]}),
    .c({\t/a/EX_fun7 [2],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b7/B9 ,\t/a/reg_writedat [7]}),
    .mi({open_n6804,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/B9 }),
    .q({open_n6819,\t/a/regfile/regfile$5$ [7]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1995|t/a/regfile/reg0_b166  (
    .a({open_n6820,_al_u1993_o}),
    .b({_al_u1985_o,\t/a/alu_B_select [1]}),
    .c({\t/a/EX_fun7 [1],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b6/B9 ,\t/a/reg_writedat [6]}),
    .mi({open_n6831,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b6/B9 }),
    .q({open_n6835,\t/a/regfile/regfile$5$ [6]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111100110000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1998|t/a/regfile/reg0_b165  (
    .a({open_n6836,_al_u1996_o}),
    .b({_al_u1985_o,\t/a/alu_B_select [1]}),
    .c({\t/a/EX_fun7 [0],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b5/B9 ,\t/a/reg_writedat [5]}),
    .mi({open_n6847,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b5/B9 }),
    .q({open_n6851,\t/a/regfile/regfile$5$ [5]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~A*~(D*~(~C*B)))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~A*~(D*~(~C*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111101110101010),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111101110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2004|t/a/regfile/reg0_b159  (
    .a({\t/a/aluin/sel1_b31/B9 ,_al_u2002_o}),
    .b({_al_u1983_o,\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [6],\t/a/reg_writedat [31]}),
    .mi({open_n6855,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [31],\t/a/aluin/sel1_b31/B9 }),
    .q({open_n6870,\t/a/regfile/regfile$4$ [31]}));  // register.v(63)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2007|t/a/id_ex/reg2_b6  (
    .c({\t/a/EX_fun7 [6],\t/a/ID_fun7 [6]}),
    .clk(clock_pad),
    .d({_al_u1983_o,\t/a/condition/n1_lutinv }),
    .mi({open_n6879,\t/a/ID_fun7 [6]}),
    .sr(rst_pad),
    .f({_al_u2007_o,\t/a/condition/sel0_b12/B1 }),
    .q({open_n6894,\t/a/EX_fun7 [6]}));  // flow_line_reg.v(139)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~B*~A*~(D*C))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111111011101110),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2008|t/a/regfile/reg0_b158  (
    .a({\t/a/aluin/sel1_b30/B9 ,_al_u2005_o}),
    .b({_al_u2007_o,\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [5],\t/a/reg_writedat [30]}),
    .mi({open_n6898,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [30],\t/a/aluin/sel1_b30/B9 }),
    .q({open_n6913,\t/a/regfile/regfile$4$ [30]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111011101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2014|t/a/regfile/reg0_b157  (
    .a({\t/a/aluin/sel1_b29/B9 ,_al_u2012_o}),
    .b({_al_u2007_o,\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [4],\t/a/reg_writedat [29]}),
    .mi({open_n6924,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [29],\t/a/aluin/sel1_b29/B9 }),
    .q({open_n6928,\t/a/regfile/regfile$4$ [29]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111011101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2017|t/a/regfile/reg0_b156  (
    .a({\t/a/aluin/sel1_b28/B9 ,_al_u2015_o}),
    .b({_al_u2007_o,\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [3],\t/a/reg_writedat [28]}),
    .mi({open_n6939,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [28],\t/a/aluin/sel1_b28/B9 }),
    .q({open_n6943,\t/a/regfile/regfile$4$ [28]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~B*~A*~(D*C))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111111011101110),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2020|t/a/regfile/reg0_b155  (
    .a({\t/a/aluin/sel1_b27/B9 ,_al_u2018_o}),
    .b({_al_u2007_o,\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [2],\t/a/reg_writedat [27]}),
    .mi({open_n6947,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [27],\t/a/aluin/sel1_b27/B9 }),
    .q({open_n6962,\t/a/regfile/regfile$4$ [27]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~B*~A*~(D*C))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111111011101110),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2023|t/a/regfile/reg0_b154  (
    .a({\t/a/aluin/sel1_b26/B9 ,_al_u2021_o}),
    .b({_al_u2007_o,\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [1],\t/a/reg_writedat [26]}),
    .mi({open_n6966,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [26],\t/a/aluin/sel1_b26/B9 }),
    .q({open_n6981,\t/a/regfile/regfile$4$ [26]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111011101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2026|t/a/regfile/reg0_b153  (
    .a({\t/a/aluin/sel1_b25/B9 ,_al_u2024_o}),
    .b({_al_u2007_o,\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_fun7 [0],\t/a/reg_writedat [25]}),
    .mi({open_n6992,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [25],\t/a/aluin/sel1_b25/B9 }),
    .q({open_n6996,\t/a/regfile/regfile$4$ [25]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("~(~B*~A*~(D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b1111111011101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2041|t/a/regfile/reg0_b148  (
    .a({\t/a/aluin/sel1_b20/B9 ,_al_u2039_o}),
    .b({_al_u2007_o,\t/a/alu_B_select [1]}),
    .c({_al_u1803_o,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/EX_rs2 [0],\t/a/reg_writedat [20]}),
    .mi({open_n7007,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [20],\t/a/aluin/sel1_b20/B9 }),
    .q({open_n7011,\t/a/regfile/regfile$4$ [20]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~D*(B@A)))"),
    //.LUT1("~(~B*~A*~(D*C))"),
    .INIT_LUT0(16'b1111000010010000),
    .INIT_LUT1(16'b1111111011101110),
    .MODE("LOGIC"))
    \_al_u2059|_al_u2445  (
    .a({\t/a/aluin/sel1_b14/B9 ,\t/a/EX_A [14]}),
    .b({_al_u2007_o,\t/a/EX_B [14]}),
    .c({_al_u1803_o,_al_u2431_o}),
    .d({\t/a/EX_fun3 [2],\t/a/EX_operation [0]}),
    .f({\t/a/EX_B [14],_al_u2445_o}));
  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("~(~B*~A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111111011101110),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2062|t/a/ex_mem/reg3_b1  (
    .a({\t/a/aluin/sel1_b13/B9 ,open_n7032}),
    .b({_al_u2007_o,open_n7033}),
    .c({_al_u1803_o,\t/a/EX_fun3 [1]}),
    .clk(clock_pad),
    .d({\t/a/EX_fun3 [1],\t/a/EX_operation [2]}),
    .mi({open_n7045,\t/a/EX_fun3 [1]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [13],_al_u2169_o}),
    .q({open_n7049,\t/a/MEM_fun3 [1]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~D*(B@A)))"),
    //.LUTF1("~(~B*~A*~(D*C))"),
    //.LUTG0("(C*~(~D*(B@A)))"),
    //.LUTG1("~(~B*~A*~(D*C))"),
    .INIT_LUTF0(16'b1111000010010000),
    .INIT_LUTF1(16'b1111111011101110),
    .INIT_LUTG0(16'b1111000010010000),
    .INIT_LUTG1(16'b1111111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2065|_al_u2465  (
    .a({\t/a/aluin/sel1_b12/B9 ,\t/a/EX_A [12]}),
    .b({_al_u2007_o,\t/a/EX_B [12]}),
    .c({_al_u1803_o,_al_u2431_o}),
    .d({\t/a/EX_fun3 [0],\t/a/EX_operation [0]}),
    .f({\t/a/EX_B [12],_al_u2465_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~D*(B@A)))"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(C*~(~D*(B@A)))"),
    //.LUTG1("~(~D*~(C*~B))"),
    .INIT_LUTF0(16'b1111000010010000),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b1111000010010000),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2068|_al_u2475  (
    .a({open_n7074,\t/a/EX_A [11]}),
    .b({_al_u1985_o,\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_fun7 [6],_al_u2431_o}),
    .d({\t/a/aluin/sel1_b11/B9 ,\t/a/EX_operation [0]}),
    .f({\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o ,_al_u2475_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("~(~D*~(C*~B))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("~(~D*~(C*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b1111111100110000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1111111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2071|t/a/regfile/reg0_b106  (
    .a({open_n7099,_al_u2069_o}),
    .b({_al_u1985_o,\t/a/alu_B_select [1]}),
    .c({\t/a/EX_fun7 [5],\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aluin/sel1_b10/B9 ,\t/a/reg_writedat [10]}),
    .mi({open_n7103,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b10/B9 }),
    .q({open_n7118,\t/a/regfile/regfile$3$ [10]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*~(D*~A*~(~0*B)))"),
    //.LUT1("~(C*~(D*~A*~(~1*B)))"),
    .INIT_LUT0(16'b0001111100001111),
    .INIT_LUT1(16'b0101111100001111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2077 (
    .a({_al_u2075_o,_al_u2075_o}),
    .b({\t/a/alu_B_select [1],\t/a/alu_B_select [1]}),
    .c({_al_u2076_o,_al_u2076_o}),
    .d({\t/a/aluin/n10_lutinv ,\t/a/aluin/n10_lutinv }),
    .mi({open_n7131,\t/a/reg_writedat [0]}),
    .fx({open_n7136,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }));
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2078|t/a/if_id/reg1_b6  (
    .a({_al_u1950_o,\t/a/if_id/n9 }),
    .b({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .c({\t/busarbitration/instruction [31],\t/busarbitration/instruction [31]}),
    .clk(clock_pad),
    .d({i_data[31],i_data[31]}),
    .sr(rst_pad),
    .f({_al_u2078_o,open_n7152}),
    .q({open_n7156,\t/a/ID_fun7 [6]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("~((C*B)*~((0*D))*~(A)+(C*B)*(0*D)*~(A)+~((C*B))*(0*D)*A+(C*B)*(0*D)*A)"),
    //.LUTF1("~((~C*~B)*~((~0*~D))*~(A)+(~C*~B)*(~0*~D)*~(A)+~((~C*~B))*(~0*~D)*A+(~C*~B)*(~0*~D)*A)"),
    //.LUTG0("~((C*B)*~((1*D))*~(A)+(C*B)*(1*D)*~(A)+~((C*B))*(1*D)*A+(C*B)*(1*D)*A)"),
    //.LUTG1("~((~C*~B)*~((~1*~D))*~(A)+(~C*~B)*(~1*~D)*~(A)+~((~C*~B))*(~1*~D)*A+(~C*~B)*(~1*~D)*A)"),
    .INIT_LUTF0(16'b1011111110111111),
    .INIT_LUTF1(16'b1111111001010100),
    .INIT_LUTG0(16'b0001010110111111),
    .INIT_LUTG1(16'b1111111011111110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2079|_al_u1944  (
    .a({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .b({\t/busarbitration/instruction [5],\t/busarbitration/instruction [5]}),
    .c({\t/busarbitration/instruction [6],\t/busarbitration/instruction [6]}),
    .d({i_data[6],i_data[6]}),
    .e({i_data[5],i_data[5]}),
    .f({\t/a/unconditional/eq1/or_xor_i0$5$_i1$5$_o_o_lutinv ,_al_u1944_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*C*~B*~A)"),
    //.LUT1("(~1*~D*C*~B*~A)"),
    .INIT_LUT0(16'b0000000000010000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2080 (
    .a({_al_u1948_o,_al_u1948_o}),
    .b({\t/instruction$2$_neg_lutinv ,\t/instruction$2$_neg_lutinv }),
    .c({\t/instruction$3$_neg_lutinv ,\t/instruction$3$_neg_lutinv }),
    .d({\t/instruction$4$_neg_lutinv ,\t/instruction$4$_neg_lutinv }),
    .mi({open_n7191,\t/a/unconditional/eq1/or_xor_i0$5$_i1$5$_o_o_lutinv }),
    .fx({open_n7196,_al_u2080_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUT1("~(~A*~(B*(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .INIT_LUT0(16'b1010111010101010),
    .INIT_LUT1(16'b1110111011101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2081 (
    .a({_al_u2078_o,_al_u2078_o}),
    .b({_al_u2080_o,_al_u2080_o}),
    .c({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .d({\t/busarbitration/instruction [30],\t/busarbitration/instruction [30]}),
    .mi({open_n7211,i_data[30]}),
    .fx({open_n7216,\t/a/IF_skip_addr [30]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUT1("~(~A*~(B*(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .INIT_LUT0(16'b1010111010101010),
    .INIT_LUT1(16'b1110111011101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2082 (
    .a({_al_u2078_o,_al_u2078_o}),
    .b({_al_u2080_o,_al_u2080_o}),
    .c({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .d({\t/busarbitration/instruction [29],\t/busarbitration/instruction [29]}),
    .mi({open_n7231,i_data[29]}),
    .fx({open_n7236,\t/a/IF_skip_addr [29]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUT1("~(~A*~(B*(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .INIT_LUT0(16'b1010111010101010),
    .INIT_LUT1(16'b1110111011101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2085 (
    .a({_al_u2078_o,_al_u2078_o}),
    .b({_al_u2080_o,_al_u2080_o}),
    .c({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .d({\t/busarbitration/instruction [26],\t/busarbitration/instruction [26]}),
    .mi({open_n7251,i_data[26]}),
    .fx({open_n7256,\t/a/IF_skip_addr [26]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(B*(D*~(0)*~(C)+D*0*~(C)+~(D)*0*C+D*0*C)))"),
    //.LUT1("~(~A*~(B*(D*~(1)*~(C)+D*1*~(C)+~(D)*1*C+D*1*C)))"),
    .INIT_LUT0(16'b1010111010101010),
    .INIT_LUT1(16'b1110111011101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2086 (
    .a({_al_u2078_o,_al_u2078_o}),
    .b({_al_u2080_o,_al_u2080_o}),
    .c({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .d({\t/busarbitration/instruction [25],\t/busarbitration/instruction [25]}),
    .mi({open_n7271,i_data[25]}),
    .fx({open_n7276,\t/a/IF_skip_addr [25]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(~C*B))"),
    //.LUTF1("~(~D*~(~C*B))"),
    //.LUTG0("~(~D*~(~C*B))"),
    //.LUTG1("~(~D*~(~C*B))"),
    .INIT_LUTF0(16'b1111111100001100),
    .INIT_LUTF1(16'b1111111100001100),
    .INIT_LUTG0(16'b1111111100001100),
    .INIT_LUTG1(16'b1111111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2087|_al_u2089  (
    .b({_al_u2080_o,_al_u2080_o}),
    .c({_al_u1956_o,_al_u1960_o}),
    .d({_al_u2078_o,_al_u2078_o}),
    .f({\t/a/IF_skip_addr [24],\t/a/IF_skip_addr [22]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~(~D*~(~C*B))"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b1111111100001100),
    .MODE("LOGIC"))
    \_al_u2088|_al_u1958  (
    .b({_al_u2080_o,\t/busarbitration/instruction [23]}),
    .c({_al_u1958_o,i_data[23]}),
    .d({_al_u2078_o,\t/busarbitration/n3 }),
    .f({\t/a/IF_skip_addr [23],_al_u1958_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~(~D*~(~C*B))"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~(~D*~(~C*B))"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b1111111100001100),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b1111111100001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2090|_al_u1965  (
    .b({_al_u2080_o,\t/busarbitration/instruction [21]}),
    .c({_al_u1965_o,i_data[21]}),
    .d({_al_u2078_o,\t/busarbitration/n3 }),
    .f({\t/a/IF_skip_addr [21],_al_u1965_o}));
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2095|t/a/if_id/reg5_b22  (
    .a({addr[22],open_n7353}),
    .b({addr[21],\t/a/MEM_aludat [22]}),
    .c({addr[20],\t/memstraddress [22]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[2],\t/busarbitration/n3 }),
    .mi({open_n7357,\t/memstraddress [22]}),
    .sr(rst_pad),
    .f({_al_u2095_o,addr[22]}),
    .q({open_n7372,\t/a/ID_memstraddr [22]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2096|t/a/if_id/reg5_b19  (
    .a({_al_u2095_o,open_n7373}),
    .b({addr[19],\t/a/MEM_aludat [19]}),
    .c({addr[18],\t/memstraddress [19]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[17],\t/busarbitration/n3 }),
    .e({addr[16],open_n7374}),
    .mi({open_n7376,\t/memstraddress [19]}),
    .sr(rst_pad),
    .f({_al_u2096_o,addr[19]}),
    .q({open_n7391,\t/a/ID_memstraddr [19]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*C*B*A)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(1*D*C*B*A)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2097|_al_u2101  (
    .a({open_n7392,_al_u2096_o}),
    .b({open_n7393,_al_u2097_o}),
    .c({addr[10],_al_u2098_o}),
    .d({addr[11],_al_u2099_o}),
    .e({open_n7396,_al_u2100_o}),
    .f({_al_u2097_o,_al_u2101_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2098|_al_u1738  (
    .c({addr[0],_al_u1737_o}),
    .d({addr[1],_al_u1735_o}),
    .f({_al_u2098_o,\t/a/risk_jump/n35_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2099|_al_u2100  (
    .c({addr[14],addr[12]}),
    .d({addr[15],addr[13]}),
    .f({_al_u2099_o,_al_u2100_o}));
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2102|t/a/if_id/reg5_b31  (
    .a({addr[5],open_n7469}),
    .b({addr[4],\t/a/MEM_aludat [31]}),
    .c({addr[31],\t/memstraddress [31]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[30],\t/busarbitration/n3 }),
    .mi({open_n7473,\t/memstraddress [31]}),
    .sr(rst_pad),
    .f({_al_u2102_o,addr[31]}),
    .q({open_n7488,\t/a/ID_memstraddr [31]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~C*B*~D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~C*B*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2103|t/a/if_id/reg5_b9  (
    .b({memwrite_cs,\t/a/MEM_aludat [9]}),
    .c({\t/a/MEM_aludat [9],\t/memstraddress [9]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[8],\t/busarbitration/n3 }),
    .mi({open_n7494,\t/memstraddress [9]}),
    .sr(rst_pad),
    .f({_al_u2103_o,addr[9]}),
    .q({open_n7509,\t/a/ID_memstraddr [9]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~C*B*A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2104|t/a/if_id/reg5_b7  (
    .a({_al_u2102_o,open_n7510}),
    .b({_al_u2103_o,\t/a/MEM_aludat [7]}),
    .c({addr[7],\t/memstraddress [7]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[6],\t/busarbitration/n3 }),
    .mi({open_n7521,\t/memstraddress [7]}),
    .sr(rst_pad),
    .f({_al_u2104_o,addr[7]}),
    .q({open_n7525,\t/a/ID_memstraddr [7]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2105|t/a/if_id/reg5_b29  (
    .a({addr[3],open_n7526}),
    .b({addr[29],\t/a/MEM_aludat [29]}),
    .c({addr[28],\t/memstraddress [29]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[27],\t/busarbitration/n3 }),
    .mi({open_n7537,\t/memstraddress [29]}),
    .sr(rst_pad),
    .f({_al_u2105_o,addr[29]}),
    .q({open_n7541,\t/a/ID_memstraddr [29]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2106|t/a/if_id/reg5_b26  (
    .b({open_n7544,\t/a/MEM_aludat [26]}),
    .c({addr[25],\t/memstraddress [26]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[26],\t/busarbitration/n3 }),
    .mi({open_n7548,\t/memstraddress [26]}),
    .sr(rst_pad),
    .f({_al_u2106_o,addr[26]}),
    .q({open_n7563,\t/a/ID_memstraddr [26]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2107|t/a/if_id/reg5_b24  (
    .b({open_n7566,\t/a/MEM_aludat [24]}),
    .c({addr[23],\t/memstraddress [24]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({addr[24],\t/busarbitration/n3 }),
    .mi({open_n7577,\t/memstraddress [24]}),
    .sr(rst_pad),
    .f({_al_u2107_o,addr[24]}),
    .q({open_n7581,\t/a/ID_memstraddr [24]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(0*D*C*B*A)"),
    //.LUT1("(1*D*C*B*A)"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2108 (
    .a({_al_u2101_o,_al_u2101_o}),
    .b({_al_u2104_o,_al_u2104_o}),
    .c({_al_u2105_o,_al_u2105_o}),
    .d({_al_u2106_o,_al_u2106_o}),
    .mi({open_n7594,_al_u2107_o}),
    .fx({open_n7599,n7}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1010100000100000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1010100000100000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2109|_al_u1954  (
    .a({open_n7602,_al_u1950_o}),
    .b({open_n7603,\t/busarbitration/n3 }),
    .c({_al_u2080_o,\t/busarbitration/instruction [26]}),
    .d({_al_u1950_o,i_data[26]}),
    .f({_al_u2109_o,\t/a/IF_skip_addr [6]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUTF0(16'b0000111100110011),
    .INIT_LUTF1(16'b0000111100110011),
    .INIT_LUTG0(16'b0000111100110011),
    .INIT_LUTG1(16'b0000111100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2111|_al_u2113  (
    .b(\t/busarbitration/instruction [19:18]),
    .c(i_data[19:18]),
    .d({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .f({_al_u2111_o,_al_u2113_o}));
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2112|t/a/if_id/reg3_b4  (
    .c({_al_u2111_o,_al_u2111_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [19],open_n7675}),
    .q({open_n7679,\t/a/ID_rs1 [4]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2114|t/a/if_id/reg3_b3  (
    .c({_al_u2113_o,_al_u2113_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [18],open_n7697}),
    .q({open_n7701,\t/a/ID_rs1 [3]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b0000111100110011),
    .MODE("LOGIC"))
    \_al_u2115|_al_u2119  (
    .b({\t/busarbitration/instruction [17],\t/busarbitration/instruction [15]}),
    .c({i_data[17],i_data[15]}),
    .d({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .f({_al_u2115_o,_al_u2119_o}));
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2116|t/a/if_id/reg3_b2  (
    .c({_al_u2115_o,_al_u2115_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [17],open_n7741}),
    .q({open_n7745,\t/a/ID_rs1 [2]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2118|t/a/if_id/reg3_b1  (
    .c({_al_u2117_o,_al_u2117_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [16],open_n7763}),
    .q({open_n7767,\t/a/ID_rs1 [1]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2120|t/a/if_id/reg3_b0  (
    .c({_al_u2119_o,_al_u2119_o}),
    .clk(clock_pad),
    .d({_al_u2109_o,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [15],open_n7785}),
    .q({open_n7789,\t/a/ID_rs1 [0]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0101010000010000),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0101010000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2121|t/a/if_id/reg0_b2  (
    .a({_al_u2109_o,\t/a/if_id/n9 }),
    .b({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .c({\t/busarbitration/instruction [14],\t/busarbitration/instruction [14]}),
    .clk(clock_pad),
    .d({i_data[14],i_data[14]}),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [14],open_n7807}),
    .q({open_n7811,\t/a/ID_fun3 [2]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0101010000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2122|t/a/if_id/reg0_b1  (
    .a({_al_u2109_o,\t/a/if_id/n9 }),
    .b({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .c({\t/busarbitration/instruction [13],\t/busarbitration/instruction [13]}),
    .clk(clock_pad),
    .d({i_data[13],i_data[13]}),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [13],open_n7825}),
    .q({open_n7829,\t/a/ID_fun3 [1]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0101010000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2123|t/a/if_id/reg0_b0  (
    .a({_al_u2109_o,\t/a/if_id/n9 }),
    .b({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .c({\t/busarbitration/instruction [12],\t/busarbitration/instruction [12]}),
    .clk(clock_pad),
    .d({i_data[12],i_data[12]}),
    .sr(rst_pad),
    .f({\t/a/IF_skip_addr [12],open_n7843}),
    .q({open_n7847,\t/a/ID_fun3 [0]}));  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"))
    \_al_u2124|_al_u596  (
    .a({\t/a/EX_fun7 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/EX_fun7 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/EX_fun7 [2],\t/a/regfile/regfile$4$ [27]}),
    .d({\t/a/EX_fun7 [3],\t/a/regfile/regfile$5$ [27]}),
    .f({_al_u2124_o,_al_u596_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(~0*D*C*B))"),
    //.LUTF1("(~D*C*~B*A)"),
    //.LUTG0("(~A*~(~1*D*C*B))"),
    //.LUTG1("(~D*C*~B*A)"),
    .INIT_LUTF0(16'b0001010101010101),
    .INIT_LUTF1(16'b0000000000100000),
    .INIT_LUTG0(16'b0101010101010101),
    .INIT_LUTG1(16'b0000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2125|_al_u2128  (
    .a({_al_u2124_o,_al_u2126_o}),
    .b({\t/a/EX_fun7 [4],\t/a/EX_operation [2]}),
    .c({\t/a/EX_fun7 [5],\t/a/aluin/n35_lutinv }),
    .d({\t/a/EX_fun7 [6],\t/a/EX_fun3 [0]}),
    .e({open_n7870,\t/a/EX_fun3 [1]}),
    .f({\t/a/aluin/n35_lutinv ,_al_u2128_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2130|_al_u2406  (
    .b({_al_u2128_o,_al_u2128_o}),
    .c({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .d({\t/a/alu/n6 [31],\t/a/alu/n6 [17]}),
    .f({_al_u2130_o,_al_u2406_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0001000011110000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b0111000011110000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2131|_al_u2436  (
    .a({open_n7917,\t/a/EX_A [15]}),
    .b({\t/a/EX_A [14],\t/a/EX_B [15]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation [1]}),
    .d({\t/a/EX_A [15],\t/a/EX_operation [2]}),
    .e({open_n7920,\t/a/EX_operation [0]}),
    .f({\t/a/alu/n156_lutinv ,_al_u2436_o}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~B))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2132|t/a/id_ex/reg7_b12  (
    .b({\t/a/EX_A [12],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [12]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [13],\t/a/aluin/sel0_b12/B0 }),
    .mi({open_n7954,\t/a/ID_memstraddr [12]}),
    .sr(rst_pad),
    .f({\t/a/alu/n158_lutinv ,\t/a/EX_A [12]}),
    .q({open_n7958,\t/a/EX_memstraddr [12]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u2133|_al_u2408  (
    .b({\t/a/alu/n158_lutinv ,\t/a/alu/n30_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n156_lutinv ,\t/a/alu/n28_lutinv }),
    .f({_al_u2133_o,_al_u2408_o}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~B))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(~D*~(C*~B))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100110000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1111111100110000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2134|t/a/id_ex/reg7_b10  (
    .b({\t/a/EX_A [10],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [10]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [11],\t/a/aluin/sel0_b10/B0 }),
    .mi({open_n7987,\t/a/ID_memstraddr [10]}),
    .sr(rst_pad),
    .f({\t/a/alu/n160_lutinv ,\t/a/EX_A [10]}),
    .q({open_n8002,\t/a/EX_memstraddr [10]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~D*(B@A)))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(C*~(~D*(B@A)))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1111000010010000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1111000010010000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2135|_al_u2505  (
    .a({open_n8003,\t/a/EX_A [8]}),
    .b({\t/a/EX_A [8],\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2431_o}),
    .d({\t/a/EX_A [9],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n162_lutinv ,_al_u2505_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0011000000111111),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u2136|_al_u2244  (
    .b({\t/a/alu/n162_lutinv ,\t/a/alu/n153_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n160_lutinv ,\t/a/alu/n151_lutinv }),
    .f({_al_u2136_o,_al_u2244_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0011111100110000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b0011111100110000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2137|_al_u2270  (
    .b({_al_u2136_o,\t/a/alu/n56_lutinv }),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2133_o,_al_u2269_o}),
    .f({_al_u2137_o,_al_u2270_o}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~B))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2138|t/a/id_ex/reg7_b7  (
    .b({\t/a/EX_A [6],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [7]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [7],\t/a/aluin/sel0_b7/B0 }),
    .mi({open_n8089,\t/a/ID_memstraddr [7]}),
    .sr(rst_pad),
    .f({\t/a/alu/n164_lutinv ,\t/a/EX_A [7]}),
    .q({open_n8093,\t/a/EX_memstraddr [7]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~B))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(~D*~(C*~B))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100110000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1111111100110000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2139|t/a/id_ex/reg7_b4  (
    .b({\t/a/EX_A [4],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [4]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [5],\t/a/aluin/sel0_b4/B0 }),
    .mi({open_n8100,\t/a/ID_memstraddr [4]}),
    .sr(rst_pad),
    .f({\t/a/alu/n166_lutinv ,\t/a/EX_A [4]}),
    .q({open_n8115,\t/a/EX_memstraddr [4]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u2140|_al_u2260  (
    .b({\t/a/alu/n166_lutinv ,_al_u2140_o}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .d({\t/a/alu/n164_lutinv ,_al_u2136_o}),
    .f({_al_u2140_o,_al_u2260_o}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~B))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2141|t/a/id_ex/reg7_b3  (
    .b({\t/a/EX_A [2],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [3]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [3],\t/a/aluin/sel0_b3/B0 }),
    .mi({open_n8151,\t/a/ID_memstraddr [3]}),
    .sr(rst_pad),
    .f({\t/a/alu/n168_lutinv ,\t/a/EX_A [3]}),
    .q({open_n8155,\t/a/EX_memstraddr [3]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u2143|_al_u2142  (
    .b({\t/a/alu/n170_lutinv ,\t/a/EX_A [0]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n168_lutinv ,\t/a/EX_A [1]}),
    .f({_al_u2143_o,\t/a/alu/n170_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2144|_al_u2384  (
    .b({_al_u2143_o,_al_u2383_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2140_o,_al_u2332_o}),
    .f({_al_u2144_o,_al_u2384_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2146|_al_u2161  (
    .c({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .d({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2146_o,_al_u2161_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2147|_al_u2313  (
    .c({_al_u2146_o,_al_u2146_o}),
    .d({_al_u2145_o,_al_u2312_o}),
    .f({_al_u2147_o,_al_u2313_o}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~B))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2148|t/a/id_ex/reg7_b22  (
    .b({\t/a/EX_A [22],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [22]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [23],\t/a/aluin/sel0_b22/B0 }),
    .mi({open_n8265,\t/a/ID_memstraddr [22]}),
    .sr(rst_pad),
    .f({\t/a/alu/n148_lutinv ,\t/a/EX_A [22]}),
    .q({open_n8269,\t/a/EX_memstraddr [22]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~B))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2149|t/a/id_ex/reg7_b21  (
    .b({\t/a/EX_A [20],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [21]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [21],\t/a/aluin/sel0_b21/B0 }),
    .mi({open_n8283,\t/a/ID_memstraddr [21]}),
    .sr(rst_pad),
    .f({\t/a/alu/n150_lutinv ,\t/a/EX_A [21]}),
    .q({open_n8287,\t/a/EX_memstraddr [21]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0011000000111111),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0011000000111111),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2150|_al_u2237  (
    .b({\t/a/alu/n150_lutinv ,\t/a/alu/n161_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n148_lutinv ,\t/a/alu/n159_lutinv }),
    .f({_al_u2150_o,_al_u2237_o}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~B))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(~D*~(C*~B))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100110000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1111111100110000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2151|t/a/id_ex/reg7_b19  (
    .b({\t/a/EX_A [18],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [19]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [19],\t/a/aluin/sel0_b19/B0 }),
    .mi({open_n8320,\t/a/ID_memstraddr [19]}),
    .sr(rst_pad),
    .f({\t/a/alu/n152_lutinv ,\t/a/EX_A [19]}),
    .q({open_n8335,\t/a/EX_memstraddr [19]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~B))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2152|t/a/id_ex/reg7_b17  (
    .b({\t/a/EX_A [16],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [17]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [17],\t/a/aluin/sel0_b17/B0 }),
    .mi({open_n8349,\t/a/ID_memstraddr [17]}),
    .sr(rst_pad),
    .f({\t/a/alu/n154_lutinv ,\t/a/EX_A [17]}),
    .q({open_n8353,\t/a/EX_memstraddr [17]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0011000000111111),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u2153|_al_u2221  (
    .b({\t/a/alu/n154_lutinv ,\t/a/alu/n152_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n152_lutinv ,\t/a/alu/n150_lutinv }),
    .f({_al_u2153_o,_al_u2221_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2154|_al_u2265  (
    .b({_al_u2153_o,_al_u2133_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2150_o,_al_u2153_o}),
    .f({_al_u2154_o,_al_u2265_o}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~B))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(~D*~(C*~B))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100110000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1111111100110000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2155|t/a/id_ex/reg7_b27  (
    .b({\t/a/EX_A [26],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [27]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [27],\t/a/aluin/sel0_b27/B0 }),
    .mi({open_n8404,\t/a/ID_memstraddr [27]}),
    .sr(rst_pad),
    .f({\t/a/alu/n144_lutinv ,\t/a/EX_A [27]}),
    .q({open_n8419,\t/a/EX_memstraddr [27]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2156|_al_u649  (
    .a({open_n8420,\t/a/ID_rs1 [0]}),
    .b({\t/a/EX_A [24],\t/a/ID_rs1 [1]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/regfile/regfile$4$ [24]}),
    .d({\t/a/EX_A [25],\t/a/regfile/regfile$5$ [24]}),
    .f({\t/a/alu/n146_lutinv ,_al_u649_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2157|_al_u2224  (
    .b({\t/a/alu/n146_lutinv ,\t/a/alu/n146_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n144_lutinv ,\t/a/alu/n148_lutinv }),
    .f({_al_u2157_o,_al_u2224_o}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~B))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(~D*~(C*~B))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100110000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1111111100110000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2158|t/a/id_ex/reg7_b28  (
    .b({\t/a/EX_A [28],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [28]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [29],\t/a/aluin/sel0_b28/B0 }),
    .mi({open_n8473,\t/a/ID_memstraddr [28]}),
    .sr(rst_pad),
    .f({\t/a/alu/n142_lutinv ,\t/a/EX_A [28]}),
    .q({open_n8488,\t/a/EX_memstraddr [28]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUT1("(~1*~(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    .INIT_LUT0(16'b1111001111110101),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2159 (
    .a({\t/a/EX_A [31],\t/a/EX_A [31]}),
    .b({\t/a/EX_A [30],\t/a/EX_A [30]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .mi({open_n8501,\t/a/EX_B [2]}),
    .fx({open_n8506,_al_u2159_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(~(D*B)*C)*~(0*A))"),
    //.LUT1("(~(~(D*B)*C)*~(1*A))"),
    .INIT_LUT0(16'b1100111100001111),
    .INIT_LUT1(16'b0100010100000101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2160 (
    .a({_al_u2157_o,_al_u2157_o}),
    .b({\t/a/alu/n142_lutinv ,\t/a/alu/n142_lutinv }),
    .c({_al_u2159_o,_al_u2159_o}),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .mi({open_n8521,\t/a/EX_B [2]}),
    .fx({open_n8526,\t/a/alu/n204_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    //.LUTG0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0101000011000000),
    .INIT_LUTG0(16'b0011000001010000),
    .INIT_LUTG1(16'b0101000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2162|_al_u2328  (
    .a({_al_u2154_o,_al_u2154_o}),
    .b({\t/a/alu/n204_lutinv ,_al_u2137_o}),
    .c({_al_u2161_o,_al_u2161_o}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2162_o,_al_u2328_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2163 (
    .a({\t/a/alu/n5 [31],\t/a/alu/n5 [31]}),
    .b({_al_u2147_o,_al_u2147_o}),
    .c({_al_u2162_o,_al_u2162_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n8565,\t/a/EX_operation [0]}),
    .fx({open_n8570,_al_u2163_o}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~B))"),
    //.LUT1("(~C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2164|t/a/id_ex/reg7_b31  (
    .b({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [31]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [31],\t/a/aluin/sel0_b31/B0 }),
    .mi({open_n8586,\t/a/ID_memstraddr [31]}),
    .sr(rst_pad),
    .f({\t/a/alu/n56_lutinv ,\t/a/EX_A [31]}),
    .q({open_n8590,\t/a/EX_memstraddr [31]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~D*C*A))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(B*~(~1*~D*C*A))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1100110001001100),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2168|_al_u2166  (
    .a({open_n8591,\t/a/alu/n56_lutinv }),
    .b({open_n8592,_al_u2165_o}),
    .c({\t/a/EX_operation [1],_al_u2161_o}),
    .d({_al_u2166_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .e({open_n8595,\t/a/EX_B [2]}),
    .f({_al_u2168_o,_al_u2166_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b1000000011100000),
    .MODE("LOGIC"))
    \_al_u2170|_al_u2165  (
    .a({\t/a/EX_A [31],\t/a/EX_A [31]}),
    .b({\t/a/EX_B [31],\t/a/EX_B [31]}),
    .c({_al_u2169_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [0],\t/a/EX_operation [2]}),
    .f({_al_u2170_o,_al_u2165_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2172|_al_u2369  (
    .b({_al_u2128_o,_al_u2128_o}),
    .c({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .d({\t/a/alu/n6 [30],\t/a/alu/n6 [20]}),
    .f({_al_u2172_o,_al_u2369_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~D*(B@A)))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1111000010010000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2173|_al_u2455  (
    .a({open_n8662,\t/a/EX_A [13]}),
    .b({\t/a/EX_A [13],\t/a/EX_B [13]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2431_o}),
    .d({\t/a/EX_A [14],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n157_lutinv ,_al_u2455_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u2175|_al_u2174  (
    .b({\t/a/alu/n159_lutinv ,\t/a/EX_A [11]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n157_lutinv ,\t/a/EX_A [12]}),
    .f({_al_u2175_o,\t/a/alu/n159_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~D*(B@A)))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111000010010000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2176|_al_u2485  (
    .a({open_n8705,\t/a/EX_A [10]}),
    .b({\t/a/EX_A [10],\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2431_o}),
    .d({\t/a/EX_A [9],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n161_lutinv ,_al_u2485_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2178|_al_u2177  (
    .b({\t/a/alu/n163_lutinv ,\t/a/EX_A [7]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n161_lutinv ,\t/a/EX_A [8]}),
    .f({_al_u2178_o,\t/a/alu/n163_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2179|_al_u2282  (
    .b({_al_u2178_o,_al_u2175_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2175_o,_al_u2194_o}),
    .f({_al_u2179_o,_al_u2282_o}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~B))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(~D*~(C*~B))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100110000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1111111100110000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2180|t/a/id_ex/reg7_b6  (
    .b({\t/a/EX_A [5],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [6]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [6],\t/a/aluin/sel0_b6/B0 }),
    .mi({open_n8784,\t/a/ID_memstraddr [6]}),
    .sr(rst_pad),
    .f({\t/a/alu/n165_lutinv ,\t/a/EX_A [6]}),
    .q({open_n8799,\t/a/EX_memstraddr [6]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(~D*(B@A)))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(~C*~(~D*(B@A)))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0000111100001001),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b0000111100001001),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2181|_al_u2546  (
    .a({open_n8800,\t/a/EX_A [4]}),
    .b({\t/a/EX_A [3],\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation [1]}),
    .d({\t/a/EX_A [4],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n167_lutinv ,_al_u2546_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2182|_al_u2277  (
    .b({\t/a/alu/n167_lutinv ,_al_u2182_o}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .d({\t/a/alu/n165_lutinv ,_al_u2178_o}),
    .f({_al_u2182_o,_al_u2277_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2183|_al_u2559  (
    .b({\t/a/EX_A [1],\t/a/EX_A [2]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_A [2],\t/a/EX_A [3]}),
    .f({\t/a/alu/n169_lutinv ,\t/a/alu/n45_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0011000000111111),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2186|_al_u2185  (
    .b({_al_u2185_o,_al_u2184_o}),
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2182_o,\t/a/alu/n169_lutinv }),
    .f({_al_u2186_o,_al_u2185_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~(~0*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(D*~C*~B*~(~1*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2188|_al_u2203  (
    .a({open_n8899,\t/a/alu/n5 [30]}),
    .b({open_n8900,_al_u2188_o}),
    .c({_al_u2146_o,_al_u2202_o}),
    .d({_al_u2187_o,_al_u2128_o}),
    .e({open_n8903,\t/a/EX_operation [0]}),
    .f({_al_u2188_o,_al_u2203_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1000000011100000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1000000011100000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2189|_al_u2363  (
    .a({open_n8924,\t/a/EX_A [21]}),
    .b({\t/a/EX_A [21],\t/a/EX_B [21]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [22],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n149_lutinv ,_al_u2363_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1000000011100000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1000000011100000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2190|_al_u2388  (
    .a({open_n8949,\t/a/EX_A [19]}),
    .b({\t/a/EX_A [19],\t/a/EX_B [19]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [20],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n151_lutinv ,_al_u2388_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0011000000111111),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u2191|_al_u2247  (
    .b({\t/a/alu/n151_lutinv ,\t/a/alu/n149_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n149_lutinv ,\t/a/alu/n147_lutinv }),
    .f({_al_u2191_o,_al_u2247_o}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~B))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(~D*~(C*~B))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111100110000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1111111100110000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2192|t/a/id_ex/reg7_b18  (
    .b({\t/a/EX_A [17],_al_u1806_o}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/EX_memstraddr [18]}),
    .clk(clock_pad),
    .d({\t/a/EX_A [18],\t/a/aluin/sel0_b18/B0 }),
    .mi({open_n9002,\t/a/ID_memstraddr [18]}),
    .sr(rst_pad),
    .f({\t/a/alu/n153_lutinv ,\t/a/EX_A [18]}),
    .q({open_n9017,\t/a/EX_memstraddr [18]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2193|_al_u2425  (
    .a({open_n9018,\t/a/EX_A [16]}),
    .b({\t/a/EX_A [15],\t/a/EX_B [16]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [16],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n155_lutinv ,_al_u2425_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u2194|_al_u2195  (
    .b({\t/a/alu/n155_lutinv ,_al_u2194_o}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .d({\t/a/alu/n153_lutinv ,_al_u2191_o}),
    .f({_al_u2194_o,_al_u2195_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2196|_al_u2308  (
    .a({open_n9061,\t/a/EX_A [25]}),
    .b({\t/a/EX_A [25],\t/a/EX_B [25]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [26],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n145_lutinv ,_al_u2308_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1000000011100000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1000000011100000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2197|_al_u2337  (
    .a({open_n9082,\t/a/EX_A [23]}),
    .b({\t/a/EX_A [23],\t/a/EX_B [23]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [24],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n147_lutinv ,_al_u2337_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0011000000111111),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u2198|_al_u2216  (
    .b({\t/a/alu/n147_lutinv ,\t/a/alu/n168_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n145_lutinv ,\t/a/alu/n166_lutinv }),
    .f({_al_u2198_o,_al_u2216_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1000000011100000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1000000011100000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2199|_al_u2274  (
    .a({open_n9129,\t/a/EX_A [27]}),
    .b({\t/a/EX_A [27],\t/a/EX_B [27]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [28],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n143_lutinv ,_al_u2274_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("((B*~(C)*~(0)+B*C*~(0)+~(B)*C*0+B*C*0)*~(A)*~(D)+(B*~(C)*~(0)+B*C*~(0)+~(B)*C*0+B*C*0)*A*~(D)+~((B*~(C)*~(0)+B*C*~(0)+~(B)*C*0+B*C*0))*A*D+(B*~(C)*~(0)+B*C*~(0)+~(B)*C*0+B*C*0)*A*D)"),
    //.LUTF1("(~C*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    //.LUTG0("((B*~(C)*~(1)+B*C*~(1)+~(B)*C*1+B*C*1)*~(A)*~(D)+(B*~(C)*~(1)+B*C*~(1)+~(B)*C*1+B*C*1)*A*~(D)+~((B*~(C)*~(1)+B*C*~(1)+~(B)*C*1+B*C*1))*A*D+(B*~(C)*~(1)+B*C*~(1)+~(B)*C*1+B*C*1)*A*D)"),
    //.LUTG1("(~C*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT_LUTF0(16'b1010101011001100),
    .INIT_LUTF1(16'b0000101000000011),
    .INIT_LUTG0(16'b1010101011110000),
    .INIT_LUTG1(16'b0000101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2201|_al_u2200  (
    .a({_al_u2198_o,\t/a/alu/n143_lutinv }),
    .b({\t/a/alu/n173_lutinv ,\t/a/EX_A [30]}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_A [29]}),
    .d({\t/a/EX_B [2],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({open_n9156,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2201_o,\t/a/alu/n173_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(C*~B*~(D*A))"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0001000000110000),
    .MODE("LOGIC"))
    \_al_u2202|_al_u2341  (
    .a({_al_u2195_o,_al_u2195_o}),
    .b({_al_u2201_o,_al_u2179_o}),
    .c({_al_u2161_o,_al_u2161_o}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2202_o,_al_u2341_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2205|_al_u2204  (
    .b({open_n9199,\t/a/EX_A [30]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n17_lutinv ,\t/a/EX_A [31]}),
    .f({\t/a/alu/n57_lutinv ,\t/a/alu/n17_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0011111100110000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2206|_al_u2287  (
    .b({open_n9226,\t/a/alu/n57_lutinv }),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({\t/a/alu/n57_lutinv ,_al_u2286_o}),
    .f({\t/a/alu/n106_lutinv ,_al_u2287_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0011111100110000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0011111100110000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2207|_al_u2347  (
    .b({open_n9249,\t/a/alu/n106_lutinv }),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n106_lutinv ,_al_u2346_o}),
    .f({\t/a/alu/n138_lutinv ,_al_u2347_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*(B@A)))"),
    //.LUTF1("(~D*~(B*~(C*A)))"),
    //.LUTG0("(D*~(~C*(B@A)))"),
    //.LUTG1("(~D*~(B*~(C*A)))"),
    .INIT_LUTF0(16'b1111100100000000),
    .INIT_LUTF1(16'b0000000010110011),
    .INIT_LUTG0(16'b1111100100000000),
    .INIT_LUTG1(16'b0000000010110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2209|_al_u2208  (
    .a({\t/a/alu/n138_lutinv ,\t/a/EX_A [30]}),
    .b({_al_u2208_o,\t/a/EX_B [30]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2209_o,_al_u2208_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1000000011100000),
    .MODE("LOGIC"))
    \_al_u2210|_al_u2234  (
    .a(\t/a/EX_A [30:29]),
    .b(\t/a/EX_B [30:29]),
    .c({_al_u2169_o,_al_u2169_o}),
    .d({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .f({_al_u2210_o,_al_u2234_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u2212|_al_u2356  (
    .b({_al_u2128_o,_al_u2128_o}),
    .c({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .d({\t/a/alu/n6 [29],\t/a/alu/n6 [21]}),
    .f({_al_u2212_o,_al_u2356_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b0011000000111111),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b0011000000111111),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2213|_al_u2214  (
    .b({\t/a/alu/n160_lutinv ,\t/a/alu/n164_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n158_lutinv ,\t/a/alu/n162_lutinv }),
    .f({_al_u2213_o,_al_u2214_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2215|_al_u2299  (
    .b({_al_u2214_o,_al_u2213_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2213_o,_al_u2222_o}),
    .f({_al_u2215_o,_al_u2299_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0011111100110000),
    .MODE("LOGIC"))
    \_al_u2218|_al_u2294  (
    .b({\t/a/alu/n202_lutinv ,_al_u2216_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2216_o,_al_u2214_o}),
    .f({_al_u2218_o,_al_u2294_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~(~0*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(D*~C*~B*~(~1*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2220|_al_u2227  (
    .a({open_n9414,\t/a/alu/n5 [29]}),
    .b({open_n9415,_al_u2220_o}),
    .c({_al_u2146_o,_al_u2226_o}),
    .d({_al_u2219_o,_al_u2128_o}),
    .e({open_n9418,\t/a/EX_operation [0]}),
    .f({_al_u2220_o,_al_u2227_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0011000000111111),
    .MODE("LOGIC"))
    \_al_u2222|_al_u2223  (
    .b({\t/a/alu/n156_lutinv ,_al_u2222_o}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .d({\t/a/alu/n154_lutinv ,_al_u2221_o}),
    .f({_al_u2222_o,_al_u2223_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(0)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(0)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*0+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*0)"),
    //.LUT1("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(1)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(1)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*1+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*1)"),
    .INIT_LUT0(16'b0011001100001111),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2225 (
    .a({_al_u2224_o,_al_u2224_o}),
    .b({\t/a/alu/n144_lutinv ,\t/a/alu/n144_lutinv }),
    .c({\t/a/alu/n142_lutinv ,\t/a/alu/n142_lutinv }),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .mi({open_n9473,\t/a/EX_B [2]}),
    .fx({open_n9478,_al_u2225_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0101000000110000),
    .INIT_LUTG0(16'b0011000001010000),
    .INIT_LUTG1(16'b0101000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2226|_al_u2354  (
    .a({_al_u2223_o,_al_u2223_o}),
    .b({_al_u2225_o,_al_u2215_o}),
    .c({_al_u2161_o,_al_u2161_o}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2226_o,_al_u2354_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(A*~((~D*B))*~(C)+A*(~D*B)*~(C)+~(A)*(~D*B)*C+A*(~D*B)*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111010100110101),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2228|_al_u2229  (
    .a({open_n9505,\t/a/alu/n18_lutinv }),
    .b({\t/a/EX_A [29],\t/a/EX_A [31]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_A [30],\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({\t/a/alu/n18_lutinv ,_al_u2229_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b0011111100110000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0011111100110000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2231|_al_u2360  (
    .b({open_n9528,\t/a/alu/n105_lutinv }),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n105_lutinv ,_al_u2359_o}),
    .f({\t/a/alu/n137_lutinv ,_al_u2360_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*(B@A)))"),
    //.LUTF1("(~D*~(B*~(C*A)))"),
    //.LUTG0("(D*~(~C*(B@A)))"),
    //.LUTG1("(~D*~(B*~(C*A)))"),
    .INIT_LUTF0(16'b1111100100000000),
    .INIT_LUTF1(16'b0000000010110011),
    .INIT_LUTG0(16'b1111100100000000),
    .INIT_LUTG1(16'b0000000010110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2233|_al_u2232  (
    .a({\t/a/alu/n137_lutinv ,\t/a/EX_A [29]}),
    .b({_al_u2232_o,\t/a/EX_B [29]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2233_o,_al_u2232_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u2236|_al_u2343  (
    .b({_al_u2128_o,_al_u2128_o}),
    .c({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .d({\t/a/alu/n6 [28],\t/a/alu/n6 [22]}),
    .f({_al_u2236_o,_al_u2343_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2238|_al_u2239  (
    .b({\t/a/alu/n165_lutinv ,_al_u2238_o}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .d({\t/a/alu/n163_lutinv ,_al_u2237_o}),
    .f({_al_u2238_o,_al_u2239_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~((~C*B))*~(D)+~A*(~C*B)*~(D)+~(~A)*(~C*B)*D+~A*(~C*B)*D)"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(~A*~((~C*B))*~(D)+~A*(~C*B)*~(D)+~(~A)*(~C*B)*D+~A*(~C*B)*D)"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1111001110101010),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b1111001110101010),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2240|_al_u2241  (
    .a({open_n9625,_al_u2240_o}),
    .b({\t/a/alu/n169_lutinv ,_al_u2184_o}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n167_lutinv ,\t/a/EX_B [2]}),
    .f({_al_u2240_o,_al_u2241_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2242|_al_u2367  (
    .a({open_n9650,_al_u2246_o}),
    .b({_al_u2241_o,_al_u2239_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,_al_u2161_o}),
    .d({_al_u2239_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2242_o,_al_u2367_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u2243|_al_u2263  (
    .c({_al_u2146_o,_al_u2146_o}),
    .d({_al_u2242_o,_al_u2262_o}),
    .f({_al_u2243_o,_al_u2263_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("~(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0011000000111111),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0011000000111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2245|_al_u2246  (
    .b({\t/a/alu/n157_lutinv ,_al_u2245_o}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .d({\t/a/alu/n155_lutinv ,_al_u2244_o}),
    .f({_al_u2245_o,_al_u2246_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(0)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(0)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*0+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*0)"),
    //.LUTF1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(1)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(1)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*1+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*1)"),
    //.LUTG1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b0101000000110000),
    .INIT_LUTG0(16'b1010101010101010),
    .INIT_LUTG1(16'b0101000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2249|_al_u2248  (
    .a({_al_u2246_o,_al_u2247_o}),
    .b({_al_u2248_o,\t/a/alu/n145_lutinv }),
    .c({_al_u2161_o,\t/a/alu/n143_lutinv }),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({open_n9723,\t/a/EX_B [2]}),
    .f({_al_u2249_o,_al_u2248_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2250 (
    .a({\t/a/alu/n5 [28],\t/a/alu/n5 [28]}),
    .b({_al_u2243_o,_al_u2243_o}),
    .c({_al_u2249_o,_al_u2249_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n9756,\t/a/EX_operation [0]}),
    .fx({open_n9761,_al_u2250_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2251|_al_u2257  (
    .a({open_n9764,\t/a/EX_A [28]}),
    .b({\t/a/EX_A [28],\t/a/EX_B [28]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [29],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n19_lutinv ,_al_u2257_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2252|_al_u2286  (
    .b({\t/a/alu/n19_lutinv ,\t/a/alu/n21_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n17_lutinv ,\t/a/alu/n19_lutinv }),
    .f({_al_u2252_o,_al_u2286_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2253|_al_u2254  (
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2252_o,\t/a/alu/n104_lutinv }),
    .f({\t/a/alu/n104_lutinv ,\t/a/alu/n136_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(B*~(C*A)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000010110011),
    .MODE("LOGIC"))
    \_al_u2256|_al_u2255  (
    .a({\t/a/alu/n136_lutinv ,\t/a/EX_A [28]}),
    .b({_al_u2255_o,\t/a/EX_B [28]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2256_o,_al_u2255_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2259|_al_u2330  (
    .b({_al_u2128_o,_al_u2128_o}),
    .c({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .d({\t/a/alu/n6 [27],\t/a/alu/n6 [23]}),
    .f({_al_u2259_o,_al_u2330_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2261|_al_u2379  (
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2143_o,\t/a/alu/n232_lutinv }),
    .f({\t/a/alu/n232_lutinv ,\t/a/alu/n264_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTG0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0011111100110000),
    .INIT_LUTG0(16'b0011000001010000),
    .INIT_LUTG1(16'b0011111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2262|_al_u2378  (
    .a({open_n9913,_al_u2265_o}),
    .b({\t/a/alu/n232_lutinv ,_al_u2260_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,_al_u2161_o}),
    .d({_al_u2260_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2262_o,_al_u2378_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2266|_al_u2264  (
    .a({_al_u2264_o,_al_u2150_o}),
    .b({_al_u2265_o,_al_u2157_o}),
    .c({_al_u2161_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .f({_al_u2266_o,_al_u2264_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2267 (
    .a({\t/a/alu/n5 [27],\t/a/alu/n5 [27]}),
    .b({_al_u2263_o,_al_u2263_o}),
    .c({_al_u2266_o,_al_u2266_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n9974,\t/a/EX_operation [0]}),
    .fx({open_n9979,_al_u2267_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u2269|_al_u2268  (
    .b({\t/a/alu/n20_lutinv ,\t/a/EX_A [27]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n18_lutinv ,\t/a/EX_A [28]}),
    .f({_al_u2269_o,\t/a/alu/n20_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u2271|_al_u2385  (
    .b({open_n10006,_al_u2270_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2270_o,_al_u2384_o}),
    .f({\t/a/alu/n135_lutinv ,_al_u2385_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(B*~(C*A)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000010110011),
    .MODE("LOGIC"))
    \_al_u2273|_al_u2272  (
    .a({\t/a/alu/n135_lutinv ,\t/a/EX_A [27]}),
    .b({_al_u2272_o,\t/a/EX_B [27]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2273_o,_al_u2272_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~C*D))"),
    //.LUTF1("(~B*~(~C*D))"),
    //.LUTG0("(~B*~(~C*D))"),
    //.LUTG1("(~B*~(~C*D))"),
    .INIT_LUTF0(16'b0011000000110011),
    .INIT_LUTF1(16'b0011000000110011),
    .INIT_LUTG0(16'b0011000000110011),
    .INIT_LUTG1(16'b0011000000110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2276|_al_u2310  (
    .b({_al_u2128_o,_al_u2128_o}),
    .c({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .d({\t/a/alu/n6 [26],\t/a/alu/n6 [24]}),
    .f({_al_u2276_o,_al_u2310_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2278|_al_u2391  (
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2185_o,\t/a/alu/n233_lutinv }),
    .f({\t/a/alu/n233_lutinv ,\t/a/alu/n265_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011111100110000),
    .MODE("LOGIC"))
    \_al_u2279|_al_u2390  (
    .a({open_n10101,_al_u2282_o}),
    .b({\t/a/alu/n233_lutinv ,_al_u2277_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,_al_u2161_o}),
    .d({_al_u2277_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2279_o,_al_u2390_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~(~0*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(D*~C*~B*~(~1*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2280|_al_u2284  (
    .a({open_n10122,\t/a/alu/n5 [26]}),
    .b({open_n10123,_al_u2280_o}),
    .c({_al_u2146_o,_al_u2283_o}),
    .d({_al_u2279_o,_al_u2128_o}),
    .e({open_n10126,\t/a/EX_operation [0]}),
    .f({_al_u2280_o,_al_u2284_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u2283|_al_u2281  (
    .a({_al_u2281_o,_al_u2198_o}),
    .b({_al_u2282_o,_al_u2191_o}),
    .c({_al_u2161_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .f({_al_u2283_o,_al_u2281_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1000000011100000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1000000011100000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2285|_al_u2291  (
    .a({open_n10167,\t/a/EX_A [26]}),
    .b({\t/a/EX_A [26],\t/a/EX_B [26]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [27],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n21_lutinv ,_al_u2291_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u2288|_al_u2397  (
    .b({open_n10194,_al_u2287_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2287_o,_al_u2396_o}),
    .f({\t/a/alu/n134_lutinv ,_al_u2397_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*(B@A)))"),
    //.LUTF1("(~D*~(B*~(C*A)))"),
    //.LUTG0("(D*~(~C*(B@A)))"),
    //.LUTG1("(~D*~(B*~(C*A)))"),
    .INIT_LUTF0(16'b1111100100000000),
    .INIT_LUTF1(16'b0000000010110011),
    .INIT_LUTG0(16'b1111100100000000),
    .INIT_LUTG1(16'b0000000010110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2290|_al_u2289  (
    .a({\t/a/alu/n134_lutinv ,\t/a/EX_A [26]}),
    .b({_al_u2289_o,\t/a/EX_B [26]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2290_o,_al_u2289_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"))
    \_al_u2295|_al_u2402  (
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n202_lutinv ,\t/a/alu/n234_lutinv }),
    .f({\t/a/alu/n234_lutinv ,\t/a/alu/n266_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTG0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0011111100110000),
    .INIT_LUTG0(16'b0011000001010000),
    .INIT_LUTG1(16'b0011111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2296|_al_u2404  (
    .a({open_n10263,_al_u2299_o}),
    .b({\t/a/alu/n234_lutinv ,_al_u2294_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,_al_u2161_o}),
    .d({_al_u2294_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2296_o,_al_u2404_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~(~0*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(D*~C*~B*~(~1*A))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2297|_al_u2301  (
    .a({open_n10288,\t/a/alu/n5 [25]}),
    .b({open_n10289,_al_u2297_o}),
    .c({_al_u2146_o,_al_u2300_o}),
    .d({_al_u2296_o,_al_u2128_o}),
    .e({open_n10292,\t/a/EX_operation [0]}),
    .f({_al_u2297_o,_al_u2301_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b0000110000001010),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u2300|_al_u2298  (
    .a({_al_u2298_o,_al_u2224_o}),
    .b({_al_u2299_o,_al_u2221_o}),
    .c({_al_u2161_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .f({_al_u2300_o,_al_u2298_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u2303|_al_u2302  (
    .b({\t/a/alu/n22_lutinv ,\t/a/EX_A [25]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n20_lutinv ,\t/a/EX_A [26]}),
    .f({_al_u2303_o,\t/a/alu/n22_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2304|_al_u2305  (
    .b({_al_u2229_o,open_n10357}),
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2303_o,_al_u2304_o}),
    .f({_al_u2304_o,\t/a/alu/n133_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(D*~(~C*(B@A)))"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1111100100000000),
    .MODE("LOGIC"))
    \_al_u2306|_al_u1344  (
    .a({\t/a/EX_A [25],\t/a/ID_rs2 [0]}),
    .b({\t/a/EX_B [25],\t/a/ID_rs2 [1]}),
    .c({\t/a/EX_operation [0],\t/a/regfile/regfile$4$ [25]}),
    .d({\t/a/EX_operation [2],\t/a/regfile/regfile$5$ [25]}),
    .f({_al_u2306_o,_al_u1344_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~D*~(B*~(C*A)))"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000010110011),
    .MODE("LOGIC"))
    \_al_u2307|_al_u2431  (
    .a({\t/a/alu/n133_lutinv ,open_n10398}),
    .b({_al_u2306_o,open_n10399}),
    .c({_al_u2161_o,\t/a/EX_operation [2]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .f({_al_u2307_o,_al_u2431_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~((~0*~D*B))*~(C)+~A*(~0*~D*B)*~(C)+~(~A)*(~0*~D*B)*C+~A*(~0*~D*B)*C)"),
    //.LUTF1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG0("~(~A*~((~1*~D*B))*~(C)+~A*(~1*~D*B)*~(C)+~(~A)*(~1*~D*B)*C+~A*(~1*~D*B)*C)"),
    //.LUTG1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUTF0(16'b1111101000111010),
    .INIT_LUTF1(16'b1100111111000000),
    .INIT_LUTG0(16'b1111101011111010),
    .INIT_LUTG1(16'b1100111111000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2311|_al_u2312  (
    .a({open_n10420,_al_u2311_o}),
    .b({_al_u2240_o,_al_u2184_o}),
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2238_o,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({open_n10423,\t/a/EX_B [2]}),
    .f({_al_u2311_o,_al_u2312_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2315|_al_u2415  (
    .a({open_n10444,_al_u2315_o}),
    .b({_al_u2237_o,_al_u2311_o}),
    .c({\t/a/EX_B [2],_al_u2161_o}),
    .d({_al_u2245_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2315_o,_al_u2415_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .INIT_LUTF0(16'b0000110000001010),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0000110000001010),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2316|_al_u2314  (
    .a({_al_u2314_o,_al_u2247_o}),
    .b({_al_u2315_o,_al_u2244_o}),
    .c({_al_u2161_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .f({_al_u2316_o,_al_u2314_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2317 (
    .a({\t/a/alu/n5 [24],\t/a/alu/n5 [24]}),
    .b({_al_u2313_o,_al_u2313_o}),
    .c({_al_u2316_o,_al_u2316_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n10501,\t/a/EX_operation [0]}),
    .fx({open_n10506,_al_u2317_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2318|_al_u2324  (
    .a({open_n10509,\t/a/EX_A [24]}),
    .b({\t/a/EX_A [24],\t/a/EX_B [24]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [25],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n23_lutinv ,_al_u2324_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2319|_al_u2345  (
    .b({\t/a/alu/n23_lutinv ,\t/a/alu/n25_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n21_lutinv ,\t/a/alu/n23_lutinv }),
    .f({_al_u2319_o,_al_u2345_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2320|_al_u2372  (
    .b({_al_u2319_o,_al_u2371_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2252_o,_al_u2319_o}),
    .f({_al_u2320_o,_al_u2372_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2321|_al_u2422  (
    .b({open_n10584,_al_u2421_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2320_o,_al_u2320_o}),
    .f({\t/a/alu/n132_lutinv ,_al_u2422_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*(B@A)))"),
    //.LUTF1("(~D*~(B*~(C*A)))"),
    //.LUTG0("(D*~(~C*(B@A)))"),
    //.LUTG1("(~D*~(B*~(C*A)))"),
    .INIT_LUTF0(16'b1111100100000000),
    .INIT_LUTF1(16'b0000000010110011),
    .INIT_LUTG0(16'b1111100100000000),
    .INIT_LUTG1(16'b0000000010110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2323|_al_u2322  (
    .a({\t/a/alu/n132_lutinv ,\t/a/EX_A [24]}),
    .b({_al_u2322_o,\t/a/EX_B [24]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2323_o,_al_u2322_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u2326|_al_u2145  (
    .b({open_n10635,_al_u2144_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2144_o,_al_u2137_o}),
    .f({\t/a/alu/n260_lutinv ,_al_u2145_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2327|_al_u2540  (
    .c({_al_u2146_o,_al_u2128_o}),
    .d({\t/a/alu/n260_lutinv ,_al_u2539_o}),
    .f({_al_u2327_o,_al_u2540_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2329 (
    .a({\t/a/alu/n5 [23],\t/a/alu/n5 [23]}),
    .b({_al_u2327_o,_al_u2327_o}),
    .c({_al_u2328_o,_al_u2328_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n10696,\t/a/EX_operation [0]}),
    .fx({open_n10701,_al_u2329_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2332|_al_u2331  (
    .b({\t/a/alu/n24_lutinv ,\t/a/EX_A [23]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n22_lutinv ,\t/a/EX_A [24]}),
    .f({_al_u2332_o,\t/a/alu/n24_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~A*~((~D*B))*~(C)+~A*(~D*B)*~(C)+~(~A)*(~D*B)*C+~A*(~D*B)*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("~(~A*~((~D*B))*~(C)+~A*(~D*B)*~(C)+~(~A)*(~D*B)*C+~A*(~D*B)*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111101000111010),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111101000111010),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2333|_al_u2334  (
    .a({open_n10730,_al_u2333_o}),
    .b({_al_u2332_o,\t/a/alu/n56_lutinv }),
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2269_o,\t/a/EX_B [2]}),
    .f({_al_u2333_o,_al_u2334_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(B*~(C*~A)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000001110011),
    .MODE("LOGIC"))
    \_al_u2336|_al_u2335  (
    .a({_al_u2334_o,\t/a/EX_A [23]}),
    .b({_al_u2335_o,\t/a/EX_B [23]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2336_o,_al_u2335_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1100111111000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1100111111000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2339|_al_u2187  (
    .b({open_n10777,_al_u2186_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2186_o,_al_u2179_o}),
    .f({\t/a/alu/n261_lutinv ,_al_u2187_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~(~0*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(D*~C*~B*~(~1*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2340|_al_u2342  (
    .a({open_n10802,\t/a/alu/n5 [22]}),
    .b({open_n10803,_al_u2340_o}),
    .c({_al_u2146_o,_al_u2341_o}),
    .d({\t/a/alu/n261_lutinv ,_al_u2128_o}),
    .e({open_n10806,\t/a/EX_operation [0]}),
    .f({_al_u2340_o,_al_u2342_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2344|_al_u2350  (
    .a({open_n10827,\t/a/EX_A [22]}),
    .b({\t/a/EX_A [22],\t/a/EX_B [22]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [23],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n25_lutinv ,_al_u2350_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2346|_al_u2396  (
    .b({_al_u2345_o,_al_u2395_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2286_o,_al_u2345_o}),
    .f({_al_u2346_o,_al_u2396_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(B*~(C*~A)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000001110011),
    .MODE("LOGIC"))
    \_al_u2349|_al_u2348  (
    .a({_al_u2347_o,\t/a/EX_A [22]}),
    .b({_al_u2348_o,\t/a/EX_B [22]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2349_o,_al_u2348_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("(~C*~D)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"))
    \_al_u2352|_al_u2219  (
    .b({open_n10892,_al_u2218_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2218_o,_al_u2215_o}),
    .f({\t/a/alu/n262_lutinv ,_al_u2219_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~(~0*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(D*~C*~B*~(~1*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2353|_al_u2355  (
    .a({open_n10913,\t/a/alu/n5 [21]}),
    .b({open_n10914,_al_u2353_o}),
    .c({_al_u2146_o,_al_u2354_o}),
    .d({\t/a/alu/n262_lutinv ,_al_u2128_o}),
    .e({open_n10917,\t/a/EX_operation [0]}),
    .f({_al_u2353_o,_al_u2355_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2358|_al_u2357  (
    .b({\t/a/alu/n26_lutinv ,\t/a/EX_A [21]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n24_lutinv ,\t/a/EX_A [22]}),
    .f({_al_u2358_o,\t/a/alu/n26_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2359|_al_u2409  (
    .b({_al_u2358_o,_al_u2408_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2303_o,_al_u2358_o}),
    .f({_al_u2359_o,_al_u2409_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*(B@A)))"),
    //.LUTF1("(~D*~(B*~(C*~A)))"),
    //.LUTG0("(D*~(~C*(B@A)))"),
    //.LUTG1("(~D*~(B*~(C*~A)))"),
    .INIT_LUTF0(16'b1111100100000000),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b1111100100000000),
    .INIT_LUTG1(16'b0000000001110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2362|_al_u2361  (
    .a({_al_u2360_o,\t/a/EX_A [21]}),
    .b({_al_u2361_o,\t/a/EX_B [21]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2362_o,_al_u2361_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2366|_al_u2365  (
    .c({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n263_lutinv ,_al_u2241_o}),
    .f({_al_u2366_o,\t/a/alu/n263_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2368 (
    .a({\t/a/alu/n5 [20],\t/a/alu/n5 [20]}),
    .b({_al_u2366_o,_al_u2366_o}),
    .c({_al_u2367_o,_al_u2367_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n11050,\t/a/EX_operation [0]}),
    .fx({open_n11055,_al_u2368_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2370|_al_u2376  (
    .a({open_n11058,\t/a/EX_A [20]}),
    .b({\t/a/EX_A [20],\t/a/EX_B [20]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [21],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n27_lutinv ,_al_u2376_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0000001111110011),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u2371|_al_u2395  (
    .b({\t/a/alu/n27_lutinv ,\t/a/alu/n29_lutinv }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n25_lutinv ,\t/a/alu/n27_lutinv }),
    .f({_al_u2371_o,_al_u2395_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*~(B*~(C*~A)))"),
    //.LUTF1("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    //.LUTG0("(~D*~(B*~(C*~A)))"),
    //.LUTG1("~(~D*~(B)*~(C)+~D*B*~(C)+~(~D)*B*C+~D*B*C)"),
    .INIT_LUTF0(16'b0000000001110011),
    .INIT_LUTF1(16'b0011111100110000),
    .INIT_LUTG0(16'b0000000001110011),
    .INIT_LUTG1(16'b0011111100110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2373|_al_u2375  (
    .a({open_n11101,_al_u2373_o}),
    .b({\t/a/alu/n104_lutinv ,_al_u2374_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,_al_u2161_o}),
    .d({_al_u2372_o,\t/a/EX_operation [1]}),
    .f({_al_u2373_o,_al_u2375_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(D*~(~C*(B@A)))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(D*~(~C*(B@A)))"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b1111100100000000),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b1111100100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2374|_al_u743  (
    .a({\t/a/EX_A [20],\t/a/ID_rs1 [0]}),
    .b({\t/a/EX_B [20],\t/a/ID_rs1 [1]}),
    .c({\t/a/EX_operation [0],\t/a/regfile/regfile$4$ [20]}),
    .d({\t/a/EX_operation [2],\t/a/regfile/regfile$5$ [20]}),
    .f({_al_u2374_o,_al_u743_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(A*~((~C*B))*~(0)+A*(~C*B)*~(0)+~(A)*(~C*B)*0+A*(~C*B)*0))"),
    //.LUTF1("(~B*~(A*~((D*C))*~(0)+A*(D*C)*~(0)+~(A)*(D*C)*0+A*(D*C)*0))"),
    //.LUTG0("(~D*(A*~((~C*B))*~(1)+A*(~C*B)*~(1)+~(A)*(~C*B)*1+A*(~C*B)*1))"),
    //.LUTG1("(~B*~(A*~((D*C))*~(1)+A*(D*C)*~(1)+~(A)*(D*C)*1+A*(D*C)*1))"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2380|_al_u2549  (
    .a({\t/a/alu/n5 [19],\t/a/alu/n5 [3]}),
    .b({_al_u2378_o,\t/a/alu/n264_lutinv }),
    .c({\t/a/alu/n264_lutinv ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation [1]}),
    .e({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .f({_al_u2380_o,\t/a/alu/mux0_b3/B1_0 }));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(~C*D))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b0011000000110011),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u2381|_al_u2293  (
    .b({\t/a/EX_operation [2],_al_u2128_o}),
    .c({_al_u2128_o,\t/a/EX_operation [0]}),
    .d({\t/a/alu/n6 [19],\t/a/alu/n6 [25]}),
    .f({_al_u2381_o,_al_u2293_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u2383|_al_u2382  (
    .b({\t/a/alu/n28_lutinv ,\t/a/EX_A [19]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n26_lutinv ,\t/a/EX_A [20]}),
    .f({_al_u2383_o,\t/a/alu/n28_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*(B@A)))"),
    //.LUTF1("(~D*~(B*~(C*~A)))"),
    //.LUTG0("(D*~(~C*(B@A)))"),
    //.LUTG1("(~D*~(B*~(C*~A)))"),
    .INIT_LUTF0(16'b1111100100000000),
    .INIT_LUTF1(16'b0000000001110011),
    .INIT_LUTG0(16'b1111100100000000),
    .INIT_LUTG1(16'b0000000001110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2387|_al_u2386  (
    .a({_al_u2385_o,\t/a/EX_A [19]}),
    .b({_al_u2386_o,\t/a/EX_B [19]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2387_o,_al_u2386_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(A*~((~C*B))*~(0)+A*(~C*B)*~(0)+~(A)*(~C*B)*0+A*(~C*B)*0))"),
    //.LUTF1("(~B*~(A*~((D*C))*~(0)+A*(D*C)*~(0)+~(A)*(D*C)*0+A*(D*C)*0))"),
    //.LUTG0("(~D*(A*~((~C*B))*~(1)+A*(~C*B)*~(1)+~(A)*(~C*B)*1+A*(~C*B)*1))"),
    //.LUTG1("(~B*~(A*~((D*C))*~(1)+A*(D*C)*~(1)+~(A)*(D*C)*1+A*(D*C)*1))"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b0001000100010001),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b0000001100110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2392|_al_u2558  (
    .a({\t/a/alu/n5 [18],\t/a/alu/n5 [2]}),
    .b({_al_u2390_o,\t/a/alu/n265_lutinv }),
    .c({\t/a/alu/n265_lutinv ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation [1]}),
    .e({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .f({_al_u2392_o,\t/a/alu/mux0_b2/B1_0 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~B*~(~C*~A)))"),
    //.LUT1("(~B*~(~C*D))"),
    .INIT_LUT0(16'b1100110100000000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"))
    \_al_u2393|_al_u2728  (
    .a({open_n11262,\t/a/alu/mux0_b6/B1_0 }),
    .b({\t/a/EX_operation [2],_al_u2526_o}),
    .c({_al_u2128_o,\t/a/EX_operation [2]}),
    .d({\t/a/alu/n6 [18],_al_u2128_o}),
    .f({_al_u2393_o,_al_u2728_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1000000011100000),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2394|_al_u2400  (
    .a({open_n11283,\t/a/EX_A [18]}),
    .b({\t/a/EX_A [18],\t/a/EX_B [18]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [19],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n29_lutinv ,_al_u2400_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(B*~(C*~A)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000001110011),
    .MODE("LOGIC"))
    \_al_u2399|_al_u2398  (
    .a({_al_u2397_o,\t/a/EX_A [18]}),
    .b({_al_u2398_o,\t/a/EX_B [18]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2399_o,_al_u2398_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~D*(A*~((~C*B))*~(0)+A*(~C*B)*~(0)+~(A)*(~C*B)*0+A*(~C*B)*0))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~D*(A*~((~C*B))*~(1)+A*(~C*B)*~(1)+~(A)*(~C*B)*1+A*(~C*B)*1))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000010101010),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000000000001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2403|_al_u2579  (
    .a({open_n11324,\t/a/alu/n5 [1]}),
    .b({open_n11325,\t/a/alu/n266_lutinv }),
    .c({_al_u2146_o,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n266_lutinv ,\t/a/EX_operation [1]}),
    .e({open_n11328,\t/a/EX_operation [0]}),
    .f({_al_u2403_o,\t/a/alu/mux0_b1/B1_0 }));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2405 (
    .a({\t/a/alu/n5 [17],\t/a/alu/n5 [17]}),
    .b({_al_u2403_o,_al_u2403_o}),
    .c({_al_u2404_o,_al_u2404_o}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n11361,\t/a/EX_operation [0]}),
    .fx({open_n11366,_al_u2405_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(C*(A*~(B)*~(D)+~(A)*B*~(D)+A*B*~(D)+A*B*D))"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1000000011100000),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1000000011100000),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2407|_al_u2413  (
    .a({open_n11369,\t/a/EX_A [17]}),
    .b({\t/a/EX_A [17],\t/a/EX_B [17]}),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,_al_u2169_o}),
    .d({\t/a/EX_A [18],\t/a/EX_operation [0]}),
    .f({\t/a/alu/n30_lutinv ,_al_u2413_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(B*~(C*~A)))"),
    //.LUT1("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    .INIT_LUT0(16'b0000000001110011),
    .INIT_LUT1(16'b1100111111000000),
    .MODE("LOGIC"))
    \_al_u2410|_al_u2412  (
    .a({open_n11394,_al_u2410_o}),
    .b({_al_u2304_o,_al_u2411_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,_al_u2161_o}),
    .d({_al_u2409_o,\t/a/EX_operation [1]}),
    .f({_al_u2410_o,_al_u2412_o}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(D*~(~C*(B@A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b1111100100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2411|t/a/id_ex/reg4_b2  (
    .a({\t/a/EX_A [17],\t/a/aluin/sel1_b17/B9 }),
    .b({\t/a/EX_B [17],_al_u2007_o}),
    .c({\t/a/EX_operation [0],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [2],\t/a/EX_rs1 [2]}),
    .mi({open_n11426,\t/a/ID_rs1 [2]}),
    .sr(rst_pad),
    .f({_al_u2411_o,\t/a/EX_B [17]}),
    .q({open_n11430,\t/a/EX_rs1 [2]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*B*A)"),
    //.LUTF1("(D*~(~C*~B*~(~0*A)))"),
    //.LUTG0("(~1*~D*~C*B*A)"),
    //.LUTG1("(D*~(~C*~B*~(~1*A)))"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b1111111000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1111110000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2417|_al_u2416  (
    .a({\t/a/alu/n5 [16],_al_u2184_o}),
    .b({_al_u2415_o,_al_u2146_o}),
    .c({_al_u2416_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2128_o,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/EX_operation [0],\t/a/EX_B [2]}),
    .f({_al_u2417_o,_al_u2416_o}));
  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~A)))"),
    //.LUT1("(~B*~(~C*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111110110000),
    .INIT_LUT1(16'b0011000000110011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2418|t/a/ex_mem/reg4_b16  (
    .a({open_n11453,_al_u2417_o}),
    .b({\t/a/EX_operation [2],_al_u2418_o}),
    .c({_al_u2128_o,_al_u2424_o}),
    .clk(clock_pad),
    .d({\t/a/alu/n6 [16],_al_u2425_o}),
    .sr(rst_pad),
    .f({_al_u2418_o,\t/a/aludat [16]}),
    .q({open_n11470,\t/a/MEM_aludat [16]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u2420|_al_u2419  (
    .b({\t/a/alu/n31_lutinv ,\t/a/EX_A [16]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n29_lutinv ,\t/a/EX_A [17]}),
    .f({_al_u2420_o,\t/a/alu/n31_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2421|_al_u2463  (
    .b({_al_u2420_o,_al_u2462_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2371_o,_al_u2420_o}),
    .f({_al_u2421_o,_al_u2463_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*(B@A)))"),
    //.LUT1("(~D*~(B*~(C*~A)))"),
    .INIT_LUT0(16'b1111100100000000),
    .INIT_LUT1(16'b0000000001110011),
    .MODE("LOGIC"))
    \_al_u2424|_al_u2423  (
    .a({_al_u2422_o,\t/a/EX_A [16]}),
    .b({_al_u2423_o,\t/a/EX_B [16]}),
    .c({_al_u2161_o,\t/a/EX_operation [0]}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [2]}),
    .f({_al_u2424_o,_al_u2423_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*~(A*~((~C*~B))*~(0)+A*(~C*~B)*~(0)+~(A)*(~C*~B)*0+A*(~C*~B)*0))"),
    //.LUT1("(~D*~(A*~((~C*~B))*~(1)+A*(~C*~B)*~(1)+~(A)*(~C*~B)*1+A*(~C*~B)*1))"),
    .INIT_LUT0(16'b0000000001010101),
    .INIT_LUT1(16'b0000000011111100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2427 (
    .a({\t/a/alu/n5 [15],\t/a/alu/n5 [15]}),
    .b({_al_u2145_o,_al_u2145_o}),
    .c({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n11551,\t/a/EX_operation [0]}),
    .fx({open_n11556,_al_u2427_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2429|_al_u2428  (
    .b({\t/a/alu/n32_lutinv ,\t/a/EX_A [15]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n30_lutinv ,\t/a/EX_A [16]}),
    .f({_al_u2429_o,\t/a/alu/n32_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2430|_al_u2473  (
    .b({_al_u2429_o,_al_u2472_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2383_o,_al_u2429_o}),
    .f({_al_u2430_o,_al_u2473_o}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(C*~(~D*(B@A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b1111000010010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2432|t/a/id_ex/reg4_b0  (
    .a({\t/a/EX_A [15],\t/a/aluin/sel1_b15/B9 }),
    .b({\t/a/EX_B [15],_al_u2007_o}),
    .c({_al_u2431_o,_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [0],\t/a/EX_rs1 [0]}),
    .mi({open_n11618,\t/a/ID_rs1 [0]}),
    .sr(rst_pad),
    .f({_al_u2432_o,\t/a/EX_B [15]}),
    .q({open_n11622,\t/a/EX_rs1 [0]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(~0*~D*C*A))"),
    //.LUTF1("(C*~(D*~(B*~(A)*~(0)+B*A*~(0)+~(B)*A*0+B*A*0)))"),
    //.LUTG0("(B*~(~1*~D*C*A))"),
    //.LUTG1("(C*~(D*~(B*~(A)*~(1)+B*A*~(1)+~(B)*A*1+B*A*1)))"),
    .INIT_LUTF0(16'b1100110001001100),
    .INIT_LUTF1(16'b1100000011110000),
    .INIT_LUTG0(16'b1100110011001100),
    .INIT_LUTG1(16'b1010000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2434|_al_u2433  (
    .a({_al_u2333_o,\t/a/alu/n56_lutinv }),
    .b({_al_u2430_o,_al_u2432_o}),
    .c({_al_u2433_o,_al_u2146_o}),
    .d({_al_u2161_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .f({_al_u2434_o,_al_u2433_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~D))"),
    //.LUT1("(~B*~(C*~D))"),
    .INIT_LUT0(16'b0011001100000011),
    .INIT_LUT1(16'b0011001100000011),
    .MODE("LOGIC"))
    \_al_u2435|_al_u2555  (
    .b({_al_u2434_o,_al_u2554_o}),
    .c({_al_u2126_o,_al_u2126_o}),
    .d({\t/a/alu/n6 [15],\t/a/alu/n6 [3]}),
    .f({_al_u2435_o,_al_u2555_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~(~D*A))"),
    //.LUT1("(C*~B*~(~D*A))"),
    .INIT_LUT0(16'b0011000000010000),
    .INIT_LUT1(16'b0011000000010000),
    .MODE("LOGIC"))
    \_al_u2438|_al_u2478  (
    .a({\t/a/alu/n5 [14],\t/a/alu/n5 [10]}),
    .b({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .c({_al_u2128_o,_al_u2128_o}),
    .d({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .f({_al_u2438_o,_al_u2478_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0001000011110000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0111000011110000),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2440|_al_u2439  (
    .a({open_n11687,\t/a/EX_A [14]}),
    .b({_al_u2439_o,\t/a/EX_B [14]}),
    .c({_al_u2126_o,\t/a/EX_operation [1]}),
    .d({\t/a/alu/n6 [14],\t/a/EX_operation [2]}),
    .e({open_n11690,\t/a/EX_operation [0]}),
    .f({_al_u2440_o,_al_u2439_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2442|_al_u2441  (
    .b({\t/a/alu/n33_lutinv ,\t/a/EX_A [14]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n31_lutinv ,\t/a/EX_A [15]}),
    .f({_al_u2442_o,\t/a/alu/n33_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2443|_al_u2483  (
    .b({_al_u2442_o,_al_u2482_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2395_o,_al_u2442_o}),
    .f({_al_u2443_o,_al_u2483_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2446|_al_u2444  (
    .a({_al_u2444_o,_al_u2346_o}),
    .b({\t/a/alu/n138_lutinv ,_al_u2443_o}),
    .c({_al_u2445_o,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2446_o,_al_u2444_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~B*~(~D*A))"),
    //.LUT1("(C*~B*~(~D*A))"),
    .INIT_LUT0(16'b0011000000010000),
    .INIT_LUT1(16'b0011000000010000),
    .MODE("LOGIC"))
    \_al_u2448|_al_u2508  (
    .a({\t/a/alu/n5 [13],\t/a/alu/n5 [7]}),
    .b({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .c({_al_u2128_o,_al_u2128_o}),
    .d({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .f({_al_u2448_o,_al_u2508_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0001000011110000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0111000011110000),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2450|_al_u2449  (
    .a({open_n11803,\t/a/EX_A [13]}),
    .b({_al_u2449_o,\t/a/EX_B [13]}),
    .c({_al_u2126_o,\t/a/EX_operation [1]}),
    .d({\t/a/alu/n6 [13],\t/a/EX_operation [2]}),
    .e({open_n11806,\t/a/EX_operation [0]}),
    .f({_al_u2450_o,_al_u2449_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u2452|_al_u2451  (
    .b({\t/a/alu/n34_lutinv ,\t/a/EX_A [13]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n32_lutinv ,\t/a/EX_A [14]}),
    .f({_al_u2452_o,\t/a/alu/n34_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b1111110000001100),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b1111110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2453|_al_u2493  (
    .b({_al_u2452_o,_al_u2492_o}),
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2408_o,_al_u2452_o}),
    .f({_al_u2453_o,_al_u2493_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2456|_al_u2454  (
    .a({_al_u2454_o,_al_u2359_o}),
    .b({\t/a/alu/n137_lutinv ,_al_u2453_o}),
    .c({_al_u2455_o,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2456_o,_al_u2454_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~(~D*A))"),
    //.LUTF1("(C*~B*~(~D*A))"),
    //.LUTG0("(C*~B*~(~D*A))"),
    //.LUTG1("(C*~B*~(~D*A))"),
    .INIT_LUTF0(16'b0011000000010000),
    .INIT_LUTF1(16'b0011000000010000),
    .INIT_LUTG0(16'b0011000000010000),
    .INIT_LUTG1(16'b0011000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2458|_al_u2498  (
    .a({\t/a/alu/n5 [12],\t/a/alu/n5 [8]}),
    .b({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .c({_al_u2128_o,_al_u2128_o}),
    .d({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .f({_al_u2458_o,_al_u2498_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUT1("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    .INIT_LUT0(16'b0001000011110000),
    .INIT_LUT1(16'b0111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2459 (
    .a({\t/a/EX_A [12],\t/a/EX_A [12]}),
    .b({\t/a/EX_B [12],\t/a/EX_B [12]}),
    .c({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n11935,\t/a/EX_operation [0]}),
    .fx({open_n11940,_al_u2459_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~D))"),
    //.LUT1("(~B*~(C*~D))"),
    .INIT_LUT0(16'b0011001100000011),
    .INIT_LUT1(16'b0011001100000011),
    .MODE("LOGIC"))
    \_al_u2460|_al_u2525  (
    .b({_al_u2459_o,_al_u2524_o}),
    .c({_al_u2126_o,_al_u2126_o}),
    .d({\t/a/alu/n6 [12],\t/a/alu/n6 [6]}),
    .f({_al_u2460_o,_al_u2525_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u2462|_al_u2461  (
    .b({\t/a/alu/n35_lutinv ,\t/a/EX_A [12]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n33_lutinv ,\t/a/EX_A [13]}),
    .f({_al_u2462_o,\t/a/alu/n35_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u2466|_al_u2464  (
    .a({_al_u2464_o,_al_u2372_o}),
    .b({\t/a/alu/n136_lutinv ,_al_u2463_o}),
    .c({_al_u2465_o,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2466_o,_al_u2464_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~B*~(~D*A))"),
    //.LUTF1("(C*~B*~(~D*A))"),
    //.LUTG0("(C*~B*~(~D*A))"),
    //.LUTG1("(C*~B*~(~D*A))"),
    .INIT_LUTF0(16'b0011000000010000),
    .INIT_LUTF1(16'b0011000000010000),
    .INIT_LUTG0(16'b0011000000010000),
    .INIT_LUTG1(16'b0011000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2468|_al_u2488  (
    .a({\t/a/alu/n5 [11],\t/a/alu/n5 [9]}),
    .b({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .c({_al_u2128_o,_al_u2128_o}),
    .d({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .f({_al_u2468_o,_al_u2488_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUT1("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    .INIT_LUT0(16'b0001000011110000),
    .INIT_LUT1(16'b0111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2469 (
    .a({\t/a/EX_A [11],\t/a/EX_A [11]}),
    .b({\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n12043,\t/a/EX_operation [0]}),
    .fx({open_n12048,_al_u2469_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~D))"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(~B*~(C*~D))"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0011001100000011),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2470|_al_u2564  (
    .b({_al_u2469_o,_al_u2563_o}),
    .c({_al_u2126_o,_al_u2126_o}),
    .d({\t/a/alu/n6 [11],\t/a/alu/n6 [2]}),
    .f({_al_u2470_o,_al_u2564_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2472|_al_u2471  (
    .b({\t/a/alu/n36_lutinv ,\t/a/EX_A [11]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n34_lutinv ,\t/a/EX_A [12]}),
    .f({_al_u2472_o,\t/a/alu/n36_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u2476|_al_u2474  (
    .a({_al_u2474_o,_al_u2384_o}),
    .b({\t/a/alu/n135_lutinv ,_al_u2473_o}),
    .c({_al_u2475_o,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2476_o,_al_u2474_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUT1("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    .INIT_LUT0(16'b0001000011110000),
    .INIT_LUT1(16'b0111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2479 (
    .a({\t/a/EX_A [10],\t/a/EX_A [10]}),
    .b({\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n12135,\t/a/EX_operation [0]}),
    .fx({open_n12140,_al_u2479_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~A*~(D*~B))"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(~C*~A*~(D*~B))"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0000010000000101),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2480|_al_u2709  (
    .a({open_n12143,_al_u2708_o}),
    .b({_al_u2479_o,\t/a/alu/n6 [10]}),
    .c({_al_u2126_o,_al_u2479_o}),
    .d({\t/a/alu/n6 [10],_al_u2126_o}),
    .f({_al_u2480_o,_al_u2709_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2482|_al_u2481  (
    .b({\t/a/alu/n37_lutinv ,\t/a/EX_A [10]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n35_lutinv ,\t/a/EX_A [11]}),
    .f({_al_u2482_o,\t/a/alu/n37_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2486|_al_u2484  (
    .a({_al_u2484_o,_al_u2396_o}),
    .b({\t/a/alu/n134_lutinv ,_al_u2483_o}),
    .c({_al_u2485_o,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2486_o,_al_u2484_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0001000011110000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0111000011110000),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2490|_al_u2489  (
    .a({open_n12218,\t/a/EX_A [9]}),
    .b({_al_u2489_o,\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o }),
    .c({_al_u2126_o,\t/a/EX_operation [1]}),
    .d({\t/a/alu/n6 [9],\t/a/EX_operation [2]}),
    .e({open_n12221,\t/a/EX_operation [0]}),
    .f({_al_u2490_o,_al_u2489_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(B)*~(C)+D*B*~(C)+~(D)*B*C+D*B*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1100111111000000),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u2492|_al_u2491  (
    .b({\t/a/alu/n38_lutinv ,\t/a/EX_A [10]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n36_lutinv ,\t/a/EX_A [9]}),
    .f({_al_u2492_o,\t/a/alu/n38_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(C*~A*~(D*B))"),
    //.LUTG0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(C*~A*~(D*B))"),
    .INIT_LUTF0(16'b0101000000110000),
    .INIT_LUTF1(16'b0001000001010000),
    .INIT_LUTG0(16'b0101000000110000),
    .INIT_LUTG1(16'b0001000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2496|_al_u2494  (
    .a({_al_u2494_o,_al_u2409_o}),
    .b({\t/a/alu/n133_lutinv ,_al_u2493_o}),
    .c({_al_u2495_o,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2496_o,_al_u2494_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUTF1("(~B*~(C*~D))"),
    //.LUTG0("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    //.LUTG1("(~B*~(C*~D))"),
    .INIT_LUTF0(16'b0001000011110000),
    .INIT_LUTF1(16'b0011001100000011),
    .INIT_LUTG0(16'b0111000011110000),
    .INIT_LUTG1(16'b0011001100000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2500|_al_u2499  (
    .a({open_n12288,\t/a/EX_A [8]}),
    .b({_al_u2499_o,\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o }),
    .c({_al_u2126_o,\t/a/EX_operation [1]}),
    .d({\t/a/alu/n6 [8],\t/a/EX_operation [2]}),
    .e({open_n12291,\t/a/EX_operation [0]}),
    .f({_al_u2500_o,_al_u2499_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u2502|_al_u2501  (
    .b({\t/a/alu/n39_lutinv ,\t/a/EX_A [8]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n37_lutinv ,\t/a/EX_A [9]}),
    .f({_al_u2502_o,\t/a/alu/n39_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2503|_al_u2544  (
    .a({open_n12334,_al_u2502_o}),
    .b({_al_u2502_o,_al_u2543_o}),
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2462_o,\t/a/EX_B [2]}),
    .f({_al_u2503_o,_al_u2544_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(C*~A*~(D*B))"),
    .INIT_LUT0(16'b0101000000110000),
    .INIT_LUT1(16'b0001000001010000),
    .MODE("LOGIC"))
    \_al_u2506|_al_u2504  (
    .a({_al_u2504_o,_al_u2421_o}),
    .b({\t/a/alu/n132_lutinv ,_al_u2503_o}),
    .c({_al_u2505_o,_al_u2161_o}),
    .d({_al_u2146_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2506_o,_al_u2504_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(D*(A*~(B)*~(0)+~(A)*B*~(0)+A*B*~(0)+A*B*0)))"),
    //.LUT1("(C*~(D*(A*~(B)*~(1)+~(A)*B*~(1)+A*B*~(1)+A*B*1)))"),
    .INIT_LUT0(16'b0001000011110000),
    .INIT_LUT1(16'b0111000011110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2509 (
    .a({\t/a/EX_A [7],\t/a/EX_A [7]}),
    .b({\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n12387,\t/a/EX_operation [0]}),
    .fx({open_n12392,_al_u2509_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2512|_al_u2511  (
    .b({\t/a/alu/n40_lutinv ,\t/a/EX_A [7]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n38_lutinv ,\t/a/EX_A [8]}),
    .f({_al_u2512_o,\t/a/alu/n40_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(C*~B*~(D*A))"),
    //.LUTG0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(C*~B*~(D*A))"),
    .INIT_LUTF0(16'b0000101000001100),
    .INIT_LUTF1(16'b0001000000110000),
    .INIT_LUTG0(16'b0000101000001100),
    .INIT_LUTG1(16'b0001000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2514|_al_u2513  (
    .a({_al_u2430_o,_al_u2472_o}),
    .b({_al_u2513_o,_al_u2512_o}),
    .c({_al_u2161_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .f({_al_u2514_o,_al_u2513_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(~D*(B@A)))"),
    //.LUTF1("(C*~A*~(D*~B))"),
    //.LUTG0("(C*~(~D*(B@A)))"),
    //.LUTG1("(C*~A*~(D*~B))"),
    .INIT_LUTF0(16'b1111000010010000),
    .INIT_LUTF1(16'b0100000001010000),
    .INIT_LUTG0(16'b1111000010010000),
    .INIT_LUTG1(16'b0100000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2516|_al_u2515  (
    .a({_al_u2514_o,\t/a/EX_A [7]}),
    .b({_al_u2334_o,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o }),
    .c({_al_u2515_o,_al_u2431_o}),
    .d({_al_u2146_o,\t/a/EX_operation [0]}),
    .f({_al_u2516_o,_al_u2515_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(A*~((~C*B))*~(0)+A*(~C*B)*~(0)+~(A)*(~C*B)*0+A*(~C*B)*0))"),
    //.LUT1("(~D*(A*~((~C*B))*~(1)+A*(~C*B)*~(1)+~(A)*(~C*B)*1+A*(~C*B)*1))"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2518 (
    .a({\t/a/alu/n5 [6],\t/a/alu/n5 [6]}),
    .b({\t/a/alu/n261_lutinv ,\t/a/alu/n261_lutinv }),
    .c({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .mi({open_n12481,\t/a/EX_operation [0]}),
    .fx({open_n12486,\t/a/alu/mux0_b6/B1_0 }));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUTF0(16'b1111110000001100),
    .INIT_LUTF1(16'b0000001111110011),
    .INIT_LUTG0(16'b1111110000001100),
    .INIT_LUTG1(16'b0000001111110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2520|_al_u2519  (
    .b({\t/a/alu/n41_lutinv ,\t/a/EX_A [6]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n39_lutinv ,\t/a/EX_A [7]}),
    .f({_al_u2520_o,\t/a/alu/n41_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*~B*~(0*A)))"),
    //.LUTF1("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG0("(C*~(D*~B*~(1*A)))"),
    //.LUTG1("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT_LUTF0(16'b1100000011110000),
    .INIT_LUTF1(16'b0000101000001100),
    .INIT_LUTG0(16'b1110000011110000),
    .INIT_LUTG1(16'b0000101000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2521|_al_u2523  (
    .a({_al_u2482_o,_al_u2443_o}),
    .b({_al_u2520_o,_al_u2521_o}),
    .c({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,_al_u2522_o}),
    .d({\t/a/EX_B [2],_al_u2161_o}),
    .e({open_n12517,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2521_o,_al_u2523_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(~(A)*~(B)*~(D)+~(A)*~(B)*D+A*~(B)*D+~(A)*B*D))"),
    //.LUT1("(C*~(~D*(B@A)))"),
    .INIT_LUT0(16'b0111000000010000),
    .INIT_LUT1(16'b1111000010010000),
    .MODE("LOGIC"))
    \_al_u2522|_al_u2526  (
    .a({\t/a/EX_A [6],\t/a/EX_A [6]}),
    .b({\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o }),
    .c({_al_u2431_o,\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .f({_al_u2522_o,_al_u2526_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(D*~(C*~B))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(D*~(C*~B))"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1100111100000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1100111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2524|_al_u2686  (
    .b({_al_u2347_o,open_n12560}),
    .c({_al_u2146_o,_al_u2161_o}),
    .d({_al_u2523_o,_al_u2187_o}),
    .f({_al_u2524_o,_al_u2686_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~D*(A*~((~C*B))*~(0)+A*(~C*B)*~(0)+~(A)*(~C*B)*0+A*(~C*B)*0))"),
    //.LUT1("(~D*(A*~((~C*B))*~(1)+A*(~C*B)*~(1)+~(A)*(~C*B)*1+A*(~C*B)*1))"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b0000000000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2528 (
    .a({\t/a/alu/n5 [5],\t/a/alu/n5 [5]}),
    .b({\t/a/alu/n262_lutinv ,\t/a/alu/n262_lutinv }),
    .c({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .mi({open_n12597,\t/a/EX_operation [0]}),
    .fx({open_n12602,\t/a/alu/mux0_b5/B1_0 }));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b0000001111110011),
    .MODE("LOGIC"))
    \_al_u2530|_al_u2529  (
    .b({\t/a/alu/n42_lutinv ,\t/a/EX_A [5]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/alu/n40_lutinv ,\t/a/EX_A [6]}),
    .f({_al_u2530_o,\t/a/alu/n42_lutinv }));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUT1("(C*~B*~(D*A))"),
    .INIT_LUT0(16'b0000101000001100),
    .INIT_LUT1(16'b0001000000110000),
    .MODE("LOGIC"))
    \_al_u2532|_al_u2531  (
    .a({_al_u2453_o,_al_u2492_o}),
    .b({_al_u2531_o,_al_u2530_o}),
    .c({_al_u2161_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .f({_al_u2532_o,_al_u2531_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~(~D*(B@A)))"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1111000010010000),
    .MODE("LOGIC"))
    \_al_u2533|_al_u418  (
    .a({\t/a/EX_A [5],\t/a/ID_rs1 [0]}),
    .b({\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ,\t/a/ID_rs1 [1]}),
    .c({_al_u2431_o,\t/a/regfile/regfile$4$ [5]}),
    .d({\t/a/EX_operation [0],\t/a/regfile/regfile$5$ [5]}),
    .f({_al_u2533_o,_al_u418_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(D*~B))"),
    //.LUT1("(~B*~(C*~D))"),
    .INIT_LUT0(16'b0100000001010000),
    .INIT_LUT1(16'b0011001100000011),
    .MODE("LOGIC"))
    \_al_u2535|_al_u2534  (
    .a({open_n12667,_al_u2532_o}),
    .b({_al_u2534_o,_al_u2360_o}),
    .c({_al_u2126_o,_al_u2533_o}),
    .d({\t/a/alu/n6 [5],_al_u2146_o}),
    .f({_al_u2535_o,_al_u2534_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*D)"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"))
    \_al_u2538|_al_u2707  (
    .c({_al_u2161_o,_al_u2161_o}),
    .d({\t/a/alu/n263_lutinv ,_al_u2279_o}),
    .f({_al_u2538_o,_al_u2707_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*(~(A)*~(B)*~(0)+~(A)*~(B)*0+A*~(B)*0+~(A)*B*0)))"),
    //.LUT1("(D*~(C*(~(A)*~(B)*~(1)+~(A)*~(B)*1+A*~(B)*1+~(A)*B*1)))"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1000111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2539 (
    .a({\t/a/EX_A [4],\t/a/EX_A [4]}),
    .b({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n12724,\t/a/EX_operation [0]}),
    .fx({open_n12729,_al_u2539_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~(~D*~(~B*~(~0*A))))"),
    //.LUT1("(C*~(~D*~(~B*~(~1*A))))"),
    .INIT_LUT0(16'b1111000000010000),
    .INIT_LUT1(16'b1111000000110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2541 (
    .a({\t/a/alu/n5 [4],\t/a/alu/n5 [4]}),
    .b({_al_u2538_o,_al_u2538_o}),
    .c({_al_u2540_o,_al_u2540_o}),
    .d({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .mi({open_n12744,\t/a/EX_operation [0]}),
    .fx({open_n12749,_al_u2541_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUT1("(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    .INIT_LUT0(16'b1111110000001100),
    .INIT_LUT1(16'b1111110000001100),
    .MODE("LOGIC"))
    \_al_u2542|_al_u2550  (
    .b(\t/a/EX_A [4:3]),
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d(\t/a/EX_A [5:4]),
    .f({\t/a/alu/n43_lutinv ,\t/a/alu/n44_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*C*~A*~(D*~B))"),
    //.LUTF1("(C*~B*~(D*A))"),
    //.LUTG0("(1*C*~A*~(D*~B))"),
    //.LUTG1("(C*~B*~(D*A))"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0001000000110000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b0001000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2545|_al_u2547  (
    .a({_al_u2463_o,_al_u2545_o}),
    .b({_al_u2544_o,_al_u2373_o}),
    .c({_al_u2161_o,_al_u2546_o}),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,_al_u2146_o}),
    .e({open_n12776,\t/a/EX_operation [2]}),
    .f({_al_u2545_o,_al_u2547_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u254|_al_u1046  (
    .c({\t/a/WB_regwritecs ,\t/a/WB_rd [0]}),
    .d({\t/a/WB_rd [4],\t/a/ID_rs2 [0]}),
    .f({_al_u254_o,_al_u1046_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(0)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(0)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*0+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*0)"),
    //.LUTF1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(1)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(1)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*1+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*1)"),
    //.LUTG1("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT_LUTF0(16'b0011001100001111),
    .INIT_LUTF1(16'b0101000000110000),
    .INIT_LUTG0(16'b1010101010101010),
    .INIT_LUTG1(16'b0101000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2552|_al_u2551  (
    .a({_al_u2473_o,_al_u2512_o}),
    .b({_al_u2551_o,\t/a/alu/n42_lutinv }),
    .c({_al_u2161_o,\t/a/alu/n44_lutinv }),
    .d({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({open_n12827,\t/a/EX_B [2]}),
    .f({_al_u2552_o,_al_u2551_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~D*(C@A)))"),
    //.LUT1("(C*~B*~(D*~A))"),
    .INIT_LUT0(16'b1100110010000100),
    .INIT_LUT1(16'b0010000000110000),
    .MODE("LOGIC"))
    \_al_u2554|_al_u2553  (
    .a({_al_u2385_o,\t/a/EX_A [3]}),
    .b({_al_u2552_o,_al_u2431_o}),
    .c({_al_u2553_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2146_o,\t/a/EX_operation [0]}),
    .f({_al_u2554_o,_al_u2553_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(0)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(0)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*0+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*0)"),
    //.LUT1("(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*~(A)*~(1)+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*~(1)+~(~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))*A*1+~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)*A*1)"),
    .INIT_LUT0(16'b0011001100001111),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2560 (
    .a({_al_u2520_o,_al_u2520_o}),
    .b({\t/a/alu/n43_lutinv ,\t/a/alu/n43_lutinv }),
    .c({\t/a/alu/n45_lutinv ,\t/a/alu/n45_lutinv }),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .mi({open_n12880,\t/a/EX_B [2]}),
    .fx({open_n12885,_al_u2560_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(~(A)*~(B)*~(D)+~(A)*~(B)*D+A*~(B)*D+~(A)*B*D))"),
    //.LUTF1("(B*~(~D*(C@A)))"),
    //.LUTG0("(C*(~(A)*~(B)*~(D)+~(A)*~(B)*D+A*~(B)*D+~(A)*B*D))"),
    //.LUTG1("(B*~(~D*(C@A)))"),
    .INIT_LUTF0(16'b0111000000010000),
    .INIT_LUTF1(16'b1100110010000100),
    .INIT_LUTG0(16'b0111000000010000),
    .INIT_LUTG1(16'b1100110010000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2561|_al_u2565  (
    .a({\t/a/EX_A [2],\t/a/EX_A [2]}),
    .b({_al_u2431_o,\t/a/EX_B [2]}),
    .c({\t/a/EX_B [2],\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .f({_al_u2561_o,_al_u2565_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(D*~(B*~(A)*~(0)+B*A*~(0)+~(B)*A*0+B*A*0)))"),
    //.LUTF1("(B*~(C*~D))"),
    //.LUTG0("(C*~(D*~(B*~(A)*~(1)+B*A*~(1)+~(B)*A*1+B*A*1)))"),
    //.LUTG1("(B*~(C*~D))"),
    .INIT_LUTF0(16'b1100000011110000),
    .INIT_LUTF1(16'b1100110000001100),
    .INIT_LUTG0(16'b1010000011110000),
    .INIT_LUTG1(16'b1100110000001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2563|_al_u2562  (
    .a({open_n12912,_al_u2483_o}),
    .b({_al_u2562_o,_al_u2560_o}),
    .c({_al_u2146_o,_al_u2561_o}),
    .d({_al_u2397_o,_al_u2161_o}),
    .e({open_n12915,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2563_o,_al_u2562_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*B*A)"),
    //.LUTF1("(~C*~B*~(~D*A))"),
    //.LUTG0("(~1*~D*~C*B*A)"),
    //.LUTG1("(~C*~B*~(~D*A))"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000001100000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000001100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2568|_al_u2567  (
    .a({\t/a/alu/n5 [0],_al_u2184_o}),
    .b({_al_u2567_o,_al_u2161_o}),
    .c({\t/a/EX_operation [1],\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_operation [0],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({open_n12938,\t/a/EX_B [2]}),
    .f({_al_u2568_o,_al_u2567_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*(~(A)*~(B)*~(0)+~(A)*~(B)*0+A*~(B)*0+~(A)*B*0))"),
    //.LUT1("(D*C*(~(A)*~(B)*~(1)+~(A)*~(B)*1+A*~(B)*1+~(A)*B*1))"),
    .INIT_LUT0(16'b0001000000000000),
    .INIT_LUT1(16'b0111000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2569 (
    .a({\t/a/EX_A [0],\t/a/EX_A [0]}),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/EX_operation [1],\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n12971,\t/a/EX_operation [0]}),
    .fx({open_n12976,_al_u2569_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000010010001100),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000010010001100),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u256|_al_u1712  (
    .a({open_n12979,\t/a/ID_rs2 [0]}),
    .b({open_n12980,\t/a/ID_rs2 [1]}),
    .c({\t/a/WB_regwritecs ,\t/a/regfile/regfile$22$ [0]}),
    .d({\t/a/WB_rd [4],\t/a/regfile/regfile$23$ [0]}),
    .f({_al_u256_o,_al_u1712_o}));
  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~(D*~A))"),
    //.LUTF1("(~C*~(~0*~(~B*~(D*~A))))"),
    //.LUTG0("(~C*~B*~(D*~A))"),
    //.LUTG1("(~C*~(~1*~(~B*~(D*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000011),
    .INIT_LUTF1(16'b0000001000000011),
    .INIT_LUTG0(16'b0000001000000011),
    .INIT_LUTG1(16'b0000111100001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2570|t/a/ex_mem/reg4_b0  (
    .a({\t/a/alu/n8 ,_al_u2570_o}),
    .b({_al_u2568_o,_al_u2571_o}),
    .c({_al_u2569_o,_al_u2577_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [1],_al_u2128_o}),
    .e({\t/a/EX_operation [2],open_n13006}),
    .sr(rst_pad),
    .f({_al_u2570_o,\t/a/aludat [0]}),
    .q({open_n13024,\t/a/MEM_aludat [0]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~D))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~B*~(C*~D))"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0011001100000011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0011001100000011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2571|_al_u2510  (
    .b({open_n13027,_al_u2509_o}),
    .c({_al_u2126_o,_al_u2126_o}),
    .d({\t/a/alu/n6 [0],\t/a/alu/n6 [7]}),
    .f({_al_u2571_o,_al_u2510_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("~(B*~(D)*~(C)+B*D*~(C)+~(B)*D*C+B*D*C)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000001111110011),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000001111110011),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2572|_al_u2543  (
    .b({open_n13054,\t/a/alu/n43_lutinv }),
    .c({\t/a/EX_B [2],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2543_o,\t/a/alu/n41_lutinv }),
    .f({_al_u2572_o,_al_u2543_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2573|_al_u2184  (
    .c({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d(\t/a/EX_A [1:0]),
    .f({_al_u2573_o,_al_u2184_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D))"),
    //.LUTF1("(D*~((~C*~B)*~(A)*~(0)+(~C*~B)*A*~(0)+~((~C*~B))*A*0+(~C*~B)*A*0))"),
    //.LUTG0("(~1*(~(~C*~B)*~(A)*~(D)+~(~C*~B)*A*~(D)+~(~(~C*~B))*A*D+~(~C*~B)*A*D))"),
    //.LUTG1("(D*~((~C*~B)*~(A)*~(1)+(~C*~B)*A*~(1)+~((~C*~B))*A*1+(~C*~B)*A*1))"),
    .INIT_LUTF0(16'b1010101011111100),
    .INIT_LUTF1(16'b1111110000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0101010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2575|_al_u2574  (
    .a({_al_u2503_o,\t/a/alu/n45_lutinv }),
    .b({_al_u2572_o,_al_u2573_o}),
    .c({_al_u2574_o,_al_u2184_o}),
    .d({_al_u2161_o,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2]}),
    .f({_al_u2575_o,_al_u2574_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(~D*(C@A)))"),
    //.LUT1("(C*~B*~(D*~A))"),
    .INIT_LUT0(16'b1100110010000100),
    .INIT_LUT1(16'b0010000000110000),
    .MODE("LOGIC"))
    \_al_u2577|_al_u2576  (
    .a({_al_u2422_o,\t/a/EX_A [0]}),
    .b({_al_u2575_o,_al_u2431_o}),
    .c({_al_u2576_o,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .d({_al_u2146_o,\t/a/EX_operation [0]}),
    .f({_al_u2577_o,_al_u2576_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(C*~D)"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2580|_al_u2230  (
    .c({\t/a/EX_B [2],\t/a/EX_B [2]}),
    .d({_al_u2530_o,_al_u2229_o}),
    .f({_al_u2580_o,\t/a/alu/n105_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTF1("(~D*~B*~(C*~A))"),
    //.LUTG0("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    //.LUTG1("(~D*~B*~(C*~A))"),
    .INIT_LUTF0(16'b0000010100000011),
    .INIT_LUTF1(16'b0000000000100011),
    .INIT_LUTG0(16'b0000010100000011),
    .INIT_LUTG1(16'b0000000000100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2582|_al_u2581  (
    .a({\t/a/alu/n44_lutinv ,\t/a/EX_A [2]}),
    .b({_al_u2581_o,\t/a/EX_A [1]}),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .d({\t/a/EX_B [2],\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({_al_u2582_o,_al_u2581_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~((~C*~B)*~(A)*~(0)+(~C*~B)*A*~(0)+~((~C*~B))*A*0+(~C*~B)*A*0))"),
    //.LUT1("(D*~((~C*~B)*~(A)*~(1)+(~C*~B)*A*~(1)+~((~C*~B))*A*1+(~C*~B)*A*1))"),
    .INIT_LUT0(16'b1111110000000000),
    .INIT_LUT1(16'b0101010100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2583 (
    .a({_al_u2493_o,_al_u2493_o}),
    .b({_al_u2580_o,_al_u2580_o}),
    .c({_al_u2582_o,_al_u2582_o}),
    .d({_al_u2161_o,_al_u2161_o}),
    .mi({open_n13213,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .fx({open_n13218,_al_u2583_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(~(A)*~(B)*~(D)+~(A)*~(B)*D+A*~(B)*D+~(A)*B*D))"),
    //.LUTF1("(B*~(~D*(C@A)))"),
    //.LUTG0("(C*(~(A)*~(B)*~(D)+~(A)*~(B)*D+A*~(B)*D+~(A)*B*D))"),
    //.LUTG1("(B*~(~D*(C@A)))"),
    .INIT_LUTF0(16'b0111000000010000),
    .INIT_LUTF1(16'b1100110010000100),
    .INIT_LUTG0(16'b0111000000010000),
    .INIT_LUTG1(16'b1100110010000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2584|_al_u2587  (
    .a({\t/a/EX_A [1],\t/a/EX_A [1]}),
    .b({_al_u2431_o,\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .c({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/EX_operation [1]}),
    .d({\t/a/EX_operation [0],\t/a/EX_operation [0]}),
    .f({_al_u2584_o,_al_u2587_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~D*~C*~A))"),
    //.LUTF1("(C*~B*~(D*~A))"),
    //.LUTG0("(~B*~(~D*~C*~A))"),
    //.LUTG1("(C*~B*~(D*~A))"),
    .INIT_LUTF0(16'b0011001100110010),
    .INIT_LUTF1(16'b0010000000110000),
    .INIT_LUTG0(16'b0011001100110010),
    .INIT_LUTG1(16'b0010000000110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2585|_al_u2586  (
    .a({_al_u2410_o,\t/a/alu/n6 [1]}),
    .b({_al_u2583_o,_al_u2585_o}),
    .c({_al_u2584_o,_al_u2128_o}),
    .d({_al_u2146_o,\t/a/EX_operation [0]}),
    .f({_al_u2585_o,_al_u2586_o}));
  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUT1("(A*~(~B*~(~D*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111001001010000),
    .INIT_LUT1(16'b1000100010001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2589|t/a/mem_wb/reg0_b6  (
    .a({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({_al_u1908_o,_al_u1908_o}),
    .c({i_data[3],\t/a/MEM_aludat [6]}),
    .clk(clock_pad),
    .d({i_data[6],i_data[6]}),
    .sr(rst_pad),
    .f({_al_u2589_o,open_n13282}),
    .q({open_n13286,\t/a/reg_writedat [6]}));  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUT1("(~A*~(~D*~C*~B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111001001010000),
    .INIT_LUT1(16'b0101010101010100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2590|t/a/mem_wb/reg0_b5  (
    .a({_al_u1908_o,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({i_data[0],_al_u1908_o}),
    .c({i_data[5],\t/a/MEM_aludat [5]}),
    .clk(clock_pad),
    .d({i_data[4],i_data[5]}),
    .sr(rst_pad),
    .f({_al_u2590_o,open_n13300}),
    .q({open_n13304,\t/a/reg_writedat [5]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(~D*C*~B*~(~0*A))"),
    //.LUT1("(~D*C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000000010000),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2591 (
    .a({\t/a/mux4_b7/B0_0 ,\t/a/mux4_b7/B0_0 }),
    .b({_al_u1904_o,_al_u1904_o}),
    .c({_al_u2589_o,_al_u2589_o}),
    .d({_al_u2590_o,_al_u2590_o}),
    .mi({open_n13317,_al_u1908_o}),
    .fx({open_n13322,_al_u2591_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~0*~D*~C*~B))"),
    //.LUT1("(A*~(~1*~D*~C*~B))"),
    .INIT_LUT0(16'b1010101010101000),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2592 (
    .a({_al_u1918_o,_al_u1918_o}),
    .b({i_data[27],i_data[27]}),
    .c({i_data[31],i_data[31]}),
    .d({i_data[29],i_data[29]}),
    .mi({open_n13337,i_data[28]}),
    .fx({open_n13342,_al_u2592_o}));
  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUTF1("(~A*~(~B*~(~D*~C)))"),
    //.LUTG0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUTG1("(~A*~(~B*~(~D*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111001001010000),
    .INIT_LUTF1(16'b0100010001000101),
    .INIT_LUTG0(16'b0111001001010000),
    .INIT_LUTG1(16'b0100010001000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2593|t/a/mem_wb/reg0_b1  (
    .a({_al_u1940_o,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({_al_u1908_o,_al_u1908_o}),
    .c({i_data[2],\t/a/MEM_aludat [1]}),
    .clk(clock_pad),
    .d({i_data[1],i_data[1]}),
    .sr(rst_pad),
    .f({_al_u2593_o,open_n13362}),
    .q({open_n13366,\t/a/reg_writedat [1]}));  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*~C))"),
    //.LUT1("(~D*C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111111101110),
    .INIT_LUT1(16'b0000000000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2594|t/a/mem_wb/reg0_b8  (
    .a({_al_u2591_o,_al_u1902_o}),
    .b({_al_u2592_o,_al_u1906_o}),
    .c({_al_u2593_o,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({_al_u1906_o,\t/a/MEM_aludat [8]}),
    .sr(rst_pad),
    .f({_al_u2594_o,open_n13380}),
    .q({open_n13384,\t/a/reg_writedat [8]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~(~C*~B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~(~C*~B))"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000011111100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2595|_al_u2890  (
    .b({i_data[14],\t/a/instr/n12 [0]}),
    .c({i_data[13],\t/memstraddress [0]}),
    .d({_al_u1903_o,_al_u2109_o}),
    .f({_al_u2595_o,_al_u2890_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u2597|_al_u1964  (
    .a({open_n13411,_al_u1950_o}),
    .b({i_data[26],\t/busarbitration/n3 }),
    .c({i_data[30],\t/busarbitration/instruction [30]}),
    .d({_al_u1918_o,i_data[30]}),
    .f({_al_u2597_o,\t/a/IF_skip_addr [10]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(~0*~D*~C*~B))"),
    //.LUT1("(A*~(~1*~D*~C*~B))"),
    .INIT_LUT0(16'b1010101010101000),
    .INIT_LUT1(16'b1010101010101010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2598 (
    .a({_al_u1918_o,_al_u1918_o}),
    .b({i_data[18],i_data[18]}),
    .c({i_data[16],i_data[16]}),
    .d({i_data[23],i_data[23]}),
    .mi({open_n13444,i_data[21]}),
    .fx({open_n13449,_al_u2598_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*A)"),
    //.LUT1("(~1*~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2599 (
    .a({_al_u2594_o,_al_u2594_o}),
    .b({_al_u2595_o,_al_u2595_o}),
    .c({_al_u2596_o,_al_u2596_o}),
    .d({_al_u2597_o,_al_u2597_o}),
    .mi({open_n13464,_al_u2598_o}),
    .fx({open_n13469,_al_u2599_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(D*~(~C*~B))"),
    .INIT_LUT0(16'b0000111100110011),
    .INIT_LUT1(16'b1111110000000000),
    .MODE("LOGIC"))
    \_al_u2600|_al_u1962  (
    .b({i_data[22],\t/busarbitration/instruction [20]}),
    .c({i_data[20],i_data[20]}),
    .d({_al_u1918_o,\t/busarbitration/n3 }),
    .f({_al_u2600_o,_al_u1962_o}));
  // PC.v(60)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~B*~A*~(C*~(~0*~D)))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~B*~A*~(C*~(~1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000100010001),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2601|t/a/instr/instr_nop_reg  (
    .a({_al_u2600_o,open_n13494}),
    .b({_al_u1917_o,_al_u2601_o}),
    .c({_al_u1918_o,_al_u2602_o}),
    .clk(clock_pad),
    .d({i_data[25],_al_u2599_o}),
    .e({i_data[24],open_n13496}),
    .sr(rst_pad),
    .f({_al_u2601_o,open_n13511}),
    .q({open_n13515,\t/instrnop }));  // PC.v(60)
  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*~C))"),
    //.LUT1("(~B*~(A*~(~D*~C)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111111101110),
    .INIT_LUT1(16'b0001000100010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2602|t/a/mem_wb/reg0_b15  (
    .a({_al_u1918_o,_al_u1917_o}),
    .b({_al_u1935_o,_al_u1935_o}),
    .c({i_data[19],\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({i_data[17],\t/a/MEM_aludat [15]}),
    .sr(rst_pad),
    .f({_al_u2602_o,open_n13529}),
    .q({open_n13533,\t/a/reg_writedat [15]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2605|_al_u1799  (
    .c({\t/a/condition/n1_lutinv ,\t/a/n9_lutinv }),
    .d({_al_u1797_o,_al_u1798_o}),
    .f({\t/a/risk_jump/n19 ,\t/a/alu_A_select [0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~0*~D*C*B))"),
    //.LUT1("(~A*~(~1*~D*C*B))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0101010101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2606 (
    .a({_al_u2604_o,_al_u2604_o}),
    .b({\t/a/risk_jump/n19 ,\t/a/risk_jump/n19 }),
    .c({\t/a/risk_jump/n42_lutinv ,\t/a/risk_jump/n42_lutinv }),
    .d({\t/a/risk_jump/n35_lutinv ,\t/a/risk_jump/n35_lutinv }),
    .mi({open_n13574,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .fx({open_n13579,_al_u2606_o}));
  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*~A)"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(~1*~D*~C*~B*~A)"),
    //.LUTG1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2608|t/a/ex_mem/reg0_b0  (
    .a({open_n13582,\t/a/EX_rd [0]}),
    .b({open_n13583,\t/a/EX_rd [1]}),
    .c({_al_u2607_o,\t/a/EX_rd [2]}),
    .clk(clock_pad),
    .d({\t/a/aluin/n11_lutinv ,\t/a/EX_rd [3]}),
    .e({open_n13585,\t/a/EX_rd [4]}),
    .mi({open_n13587,\t/a/EX_rd [0]}),
    .sr(rst_pad),
    .f({_al_u2608_o,_al_u2607_o}),
    .q({open_n13602,\t/a/MEM_rd [0]}));  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2610|_al_u2710  (
    .b({open_n13605,_al_u2610_o}),
    .c({_al_u2604_o,\t/a/ID_read_dat2 [10]}),
    .d({_al_u2609_o,_al_u2606_o}),
    .f({_al_u2610_o,_al_u2710_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2612|t/a/regfile/reg0_b127  (
    .a({\t/a/aludat [31],_al_u2606_o}),
    .b({_al_u2611_o,_al_u2610_o}),
    .c({_al_u2606_o,\t/a/MEM_aludat [31]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o,\t/a/reg_writedat [31]}),
    .e({\t/a/ID_read_dat2 [31],open_n13630}),
    .mi({open_n13632,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [31],_al_u2611_o}),
    .q({open_n13647,\t/a/regfile/regfile$3$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(~0*~D*C*B))"),
    //.LUT1("(~A*~(~1*~D*C*B))"),
    .INIT_LUT0(16'b0101010100010101),
    .INIT_LUT1(16'b0101010101010101),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2614 (
    .a({_al_u2613_o,_al_u2613_o}),
    .b({\t/a/risk_jump/n19 ,\t/a/risk_jump/n19 }),
    .c({\t/a/risk_jump/n24_lutinv ,\t/a/risk_jump/n24_lutinv }),
    .d({\t/a/risk_jump/n11_lutinv ,\t/a/risk_jump/n11_lutinv }),
    .mi({open_n13660,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .fx({open_n13665,_al_u2614_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(~C*~D)"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(~C*~D)"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b0000000000001111),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b0000000000001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2616|_al_u2692  (
    .b({open_n13670,_al_u2616_o}),
    .c({_al_u2613_o,\t/a/ID_read_dat1 [14]}),
    .d({_al_u2615_o,_al_u2614_o}),
    .f({_al_u2616_o,_al_u2692_o}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2618|t/a/id_ex/reg8_b31  (
    .a({\t/a/aludat [31],_al_u333_o}),
    .b({_al_u2617_o,_al_u490_o}),
    .c({_al_u2614_o,_al_u500_o}),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [31]}),
    .e({\t/a/ID_read_dat1 [31],open_n13696}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [31],\t/a/ID_read_dat1 [31]}),
    .q({open_n13714,\t/a/EX_regdat1 [31]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2622 (
    .a({\t/a/aludat [30],\t/a/aludat [30]}),
    .b({_al_u2621_o,_al_u2621_o}),
    .c({_al_u2614_o,_al_u2614_o}),
    .d({_al_u2616_o,_al_u2616_o}),
    .mi({open_n13727,\t/a/ID_read_dat1 [30]}),
    .fx({open_n13732,\t/a/ID_jump_regdat1 [30]}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2626|t/a/id_ex/reg8_b29  (
    .a({\t/a/aludat [29],_al_u333_o}),
    .b({_al_u2625_o,_al_u553_o}),
    .c({_al_u2614_o,_al_u563_o}),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [29]}),
    .e({\t/a/ID_read_dat1 [29],open_n13736}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [29],\t/a/ID_read_dat1 [29]}),
    .q({open_n13754,\t/a/EX_regdat1 [29]}));  // flow_line_reg.v(139)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2628|t/a/regfile/reg0_b124  (
    .a({\t/a/aludat [28],_al_u2606_o}),
    .b({_al_u2627_o,_al_u2610_o}),
    .c({_al_u2606_o,\t/a/MEM_aludat [28]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o,\t/a/reg_writedat [28]}),
    .e({\t/a/ID_read_dat2 [28],open_n13755}),
    .mi({open_n13757,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [28],_al_u2627_o}),
    .q({open_n13772,\t/a/regfile/regfile$3$ [28]}));  // register.v(63)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2630|t/a/id_ex/reg8_b28  (
    .a({\t/a/aludat [28],_al_u333_o}),
    .b({_al_u2629_o,_al_u574_o}),
    .c({_al_u2614_o,_al_u584_o}),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [28]}),
    .e({\t/a/ID_read_dat1 [28],open_n13774}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [28],\t/a/ID_read_dat1 [28]}),
    .q({open_n13792,\t/a/EX_regdat1 [28]}));  // flow_line_reg.v(139)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2632|t/a/regfile/reg0_b123  (
    .a({\t/a/aludat [27],_al_u2606_o}),
    .b({_al_u2631_o,_al_u2610_o}),
    .c({_al_u2606_o,\t/a/MEM_aludat [27]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o,\t/a/reg_writedat [27]}),
    .e({\t/a/ID_read_dat2 [27],open_n13793}),
    .mi({open_n13795,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [27],_al_u2631_o}),
    .q({open_n13810,\t/a/regfile/regfile$3$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2634 (
    .a({\t/a/aludat [27],\t/a/aludat [27]}),
    .b({_al_u2633_o,_al_u2633_o}),
    .c({_al_u2614_o,_al_u2614_o}),
    .d({_al_u2616_o,_al_u2616_o}),
    .mi({open_n13823,\t/a/ID_read_dat1 [27]}),
    .fx({open_n13828,\t/a/ID_jump_regdat1 [27]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2638 (
    .a({\t/a/aludat [26],\t/a/aludat [26]}),
    .b({_al_u2637_o,_al_u2637_o}),
    .c({_al_u2614_o,_al_u2614_o}),
    .d({_al_u2616_o,_al_u2616_o}),
    .mi({open_n13843,\t/a/ID_read_dat1 [26]}),
    .fx({open_n13848,\t/a/ID_jump_regdat1 [26]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2640 (
    .a({\t/a/aludat [25],\t/a/aludat [25]}),
    .b({_al_u2639_o,_al_u2639_o}),
    .c({_al_u2606_o,_al_u2606_o}),
    .d({_al_u2610_o,_al_u2610_o}),
    .mi({open_n13863,\t/a/ID_read_dat2 [25]}),
    .fx({open_n13868,\t/a/ID_jump_regdat2 [25]}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2642|t/a/id_ex/reg8_b25  (
    .a({\t/a/aludat [25],_al_u333_o}),
    .b({_al_u2641_o,_al_u637_o}),
    .c({_al_u2614_o,_al_u647_o}),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [25]}),
    .e({\t/a/ID_read_dat1 [25],open_n13872}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [25],\t/a/ID_read_dat1 [25]}),
    .q({open_n13890,\t/a/EX_regdat1 [25]}));  // flow_line_reg.v(139)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2644|t/a/regfile/reg0_b120  (
    .a({\t/a/aludat [24],_al_u2606_o}),
    .b({_al_u2643_o,_al_u2610_o}),
    .c({_al_u2606_o,\t/a/MEM_aludat [24]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o,\t/a/reg_writedat [24]}),
    .e({\t/a/ID_read_dat2 [24],open_n13891}),
    .mi({open_n13893,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [24],_al_u2643_o}),
    .q({open_n13908,\t/a/regfile/regfile$3$ [24]}));  // register.v(63)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2646|t/a/id_ex/reg8_b24  (
    .a({\t/a/aludat [24],_al_u333_o}),
    .b({_al_u2645_o,_al_u658_o}),
    .c({_al_u2614_o,_al_u668_o}),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [24]}),
    .e({\t/a/ID_read_dat1 [24],open_n13910}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [24],\t/a/ID_read_dat1 [24]}),
    .q({open_n13928,\t/a/EX_regdat1 [24]}));  // flow_line_reg.v(139)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2648|t/a/regfile/reg0_b119  (
    .a({\t/a/aludat [23],_al_u2606_o}),
    .b({_al_u2647_o,_al_u2610_o}),
    .c({_al_u2606_o,\t/a/MEM_aludat [23]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o,\t/a/reg_writedat [23]}),
    .e({\t/a/ID_read_dat2 [23],open_n13929}),
    .mi({open_n13931,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [23],_al_u2647_o}),
    .q({open_n13946,\t/a/regfile/regfile$3$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2652|_al_u2654  (
    .a({\t/a/aludat [22],\t/a/aludat [22]}),
    .b({_al_u2651_o,_al_u2653_o}),
    .c({_al_u2606_o,_al_u2614_o}),
    .d({_al_u2610_o,_al_u2616_o}),
    .e({\t/a/ID_read_dat2 [22],\t/a/ID_read_dat1 [22]}),
    .f({\t/a/ID_jump_regdat2 [22],\t/a/ID_jump_regdat1 [22]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2656 (
    .a({\t/a/aludat [21],\t/a/aludat [21]}),
    .b({_al_u2655_o,_al_u2655_o}),
    .c({_al_u2606_o,_al_u2606_o}),
    .d({_al_u2610_o,_al_u2610_o}),
    .mi({open_n13981,\t/a/ID_read_dat2 [21]}),
    .fx({open_n13986,\t/a/ID_jump_regdat2 [21]}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2658|t/a/id_ex/reg8_b21  (
    .a({\t/a/aludat [21],_al_u333_o}),
    .b({_al_u2657_o,_al_u721_o}),
    .c({_al_u2614_o,_al_u731_o}),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [21]}),
    .e({\t/a/ID_read_dat1 [21],open_n13990}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [21],\t/a/ID_read_dat1 [21]}),
    .q({open_n14008,\t/a/EX_regdat1 [21]}));  // flow_line_reg.v(139)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2660|t/a/regfile/reg0_b116  (
    .a({\t/a/aludat [20],_al_u2606_o}),
    .b({_al_u2659_o,_al_u2610_o}),
    .c({_al_u2606_o,\t/a/MEM_aludat [20]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o,\t/a/reg_writedat [20]}),
    .e({\t/a/ID_read_dat2 [20],open_n14009}),
    .mi({open_n14011,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [20],_al_u2659_o}),
    .q({open_n14026,\t/a/regfile/regfile$3$ [20]}));  // register.v(63)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2662|t/a/id_ex/reg8_b20  (
    .a({\t/a/aludat [20],_al_u333_o}),
    .b({_al_u2661_o,_al_u742_o}),
    .c({_al_u2614_o,_al_u752_o}),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [20]}),
    .e({\t/a/ID_read_dat1 [20],open_n14028}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [20],\t/a/ID_read_dat1 [20]}),
    .q({open_n14046,\t/a/EX_regdat1 [20]}));  // flow_line_reg.v(139)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2664|t/a/regfile/reg0_b115  (
    .a({\t/a/aludat [19],_al_u2606_o}),
    .b({_al_u2663_o,_al_u2610_o}),
    .c({_al_u2606_o,\t/a/MEM_aludat [19]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o,\t/a/reg_writedat [19]}),
    .e({\t/a/ID_read_dat2 [19],open_n14047}),
    .mi({open_n14049,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [19],_al_u2663_o}),
    .q({open_n14064,\t/a/regfile/regfile$3$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2666 (
    .a({\t/a/aludat [19],\t/a/aludat [19]}),
    .b({_al_u2665_o,_al_u2665_o}),
    .c({_al_u2614_o,_al_u2614_o}),
    .d({_al_u2616_o,_al_u2616_o}),
    .mi({open_n14077,\t/a/ID_read_dat1 [19]}),
    .fx({open_n14082,\t/a/ID_jump_regdat1 [19]}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2670|t/a/id_ex/reg8_b18  (
    .a({\t/a/aludat [18],_al_u333_o}),
    .b({_al_u2669_o,_al_u805_o}),
    .c({_al_u2614_o,_al_u815_o}),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [18]}),
    .e({\t/a/ID_read_dat1 [18],open_n14086}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [18],\t/a/ID_read_dat1 [18]}),
    .q({open_n14104,\t/a/EX_regdat1 [18]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2674|t/a/id_ex/reg8_b17  (
    .a({\t/a/aludat [17],_al_u333_o}),
    .b({_al_u2673_o,_al_u826_o}),
    .c({_al_u2614_o,_al_u836_o}),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [17]}),
    .e({\t/a/ID_read_dat1 [17],open_n14106}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [17],\t/a/ID_read_dat1 [17]}),
    .q({open_n14124,\t/a/EX_regdat1 [17]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2676 (
    .a({\t/a/aludat [16],\t/a/aludat [16]}),
    .b({_al_u2675_o,_al_u2675_o}),
    .c({_al_u2606_o,_al_u2606_o}),
    .d({_al_u2610_o,_al_u2610_o}),
    .mi({open_n14137,\t/a/ID_read_dat2 [16]}),
    .fx({open_n14142,\t/a/ID_jump_regdat2 [16]}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2678|t/a/regfile/reg0_b1008  (
    .a({\t/a/aludat [16],_al_u2614_o}),
    .b({_al_u2677_o,_al_u2616_o}),
    .c({_al_u2614_o,\t/a/MEM_aludat [16]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [16]}),
    .e({\t/a/ID_read_dat1 [16],open_n14145}),
    .mi({open_n14147,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [16],_al_u2677_o}),
    .q({open_n14162,\t/a/regfile/regfile$31$ [16]}));  // register.v(63)
  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(D*~(~C*~A)))"),
    //.LUTF1("(C*~(~B*~D))"),
    //.LUTG0("(B*~(D*~(~C*~A)))"),
    //.LUTG1("(C*~(~B*~D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010011001100),
    .INIT_LUTF1(16'b1111000011000000),
    .INIT_LUTG0(16'b0000010011001100),
    .INIT_LUTG1(16'b1111000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2679|t/a/ex_mem/reg4_b15  (
    .a({open_n14163,_al_u2427_o}),
    .b({_al_u2436_o,_al_u2435_o}),
    .c({_al_u2128_o,_al_u2436_o}),
    .clk(clock_pad),
    .d({_al_u2427_o,_al_u2128_o}),
    .sr(rst_pad),
    .f({_al_u2679_o,open_n14181}),
    .q({open_n14185,\t/a/MEM_aludat [15]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u2680|_al_u2748  (
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/ID_read_dat2 [15],\t/a/ID_read_dat2 [3]}),
    .d({_al_u2606_o,_al_u2606_o}),
    .f({_al_u2680_o,_al_u2748_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(B*~A))))"),
    .INIT_LUT0(16'b1111111101000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2682 (
    .a({_al_u2679_o,_al_u2679_o}),
    .b({_al_u2435_o,_al_u2435_o}),
    .c({_al_u2680_o,_al_u2680_o}),
    .d({_al_u2681_o,_al_u2681_o}),
    .mi({open_n14220,_al_u2610_o}),
    .fx({open_n14225,\t/a/ID_jump_regdat2 [15]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~(~C*B))"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("(D*~(~C*B))"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b1111001100000000),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b1111001100000000),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2683|_al_u2713  (
    .b({_al_u2616_o,_al_u2616_o}),
    .c({\t/a/ID_read_dat1 [15],\t/a/ID_read_dat1 [10]}),
    .d({_al_u2614_o,_al_u2614_o}),
    .f({_al_u2683_o,_al_u2713_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~D*~(C*~(~1*~(B*~A))))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1111111101000000),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2685|t/a/regfile/reg0_b1007  (
    .a({_al_u2679_o,_al_u2614_o}),
    .b({_al_u2435_o,_al_u2616_o}),
    .c({_al_u2683_o,\t/a/MEM_aludat [15]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2684_o,\t/a/reg_writedat [15]}),
    .e({_al_u2616_o,open_n14254}),
    .mi({open_n14256,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [15],_al_u2684_o}),
    .q({open_n14271,\t/a/regfile/regfile$31$ [15]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(D*~C*~B*~(~0*A))"),
    //.LUTF1("(~C*~A*~(D*~B))"),
    //.LUTG0("(D*~C*~B*~(~1*A))"),
    //.LUTG1("(~C*~A*~(D*~B))"),
    .INIT_LUTF0(16'b0000000100000000),
    .INIT_LUTF1(16'b0000010000000101),
    .INIT_LUTG0(16'b0000001100000000),
    .INIT_LUTG1(16'b0000010000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2688|_al_u2687  (
    .a({_al_u2687_o,\t/a/alu/n5 [14]}),
    .b({\t/a/alu/n6 [14],_al_u2686_o}),
    .c({_al_u2439_o,\t/a/EX_operation [2]}),
    .d({_al_u2126_o,_al_u2128_o}),
    .e({open_n14274,\t/a/EX_operation [0]}),
    .f({_al_u2688_o,_al_u2687_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(~C*B))"),
    //.LUT1("(D*~(~C*B))"),
    .INIT_LUT0(16'b1111001100000000),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"))
    \_al_u2690|_al_u2729  (
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/ID_read_dat2 [14],\t/a/ID_read_dat2 [6]}),
    .d({_al_u2606_o,_al_u2606_o}),
    .f({_al_u2690_o,_al_u2729_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(~0*~(~B*A))))"),
    //.LUTF1("~(~C*~(D*~(~0*~(~B*A))))"),
    //.LUTG0("~(~D*~(C*~(~1*~(~B*A))))"),
    //.LUTG1("~(~C*~(D*~(~1*~(~B*A))))"),
    .INIT_LUTF0(16'b1111111100100000),
    .INIT_LUTF1(16'b1111001011110000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2691|_al_u2694  (
    .a({_al_u2688_o,_al_u2688_o}),
    .b({_al_u2446_o,_al_u2446_o}),
    .c({_al_u2689_o,_al_u2692_o}),
    .d({_al_u2690_o,_al_u2693_o}),
    .e({_al_u2610_o,_al_u2616_o}),
    .f({\t/a/ID_jump_regdat2 [14],\t/a/ID_jump_regdat1 [14]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2696 (
    .a({\t/a/aludat [13],\t/a/aludat [13]}),
    .b({_al_u2695_o,_al_u2695_o}),
    .c({_al_u2606_o,_al_u2606_o}),
    .d({_al_u2610_o,_al_u2610_o}),
    .mi({open_n14351,\t/a/ID_read_dat2 [13]}),
    .fx({open_n14356,\t/a/ID_jump_regdat2 [13]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2698 (
    .a({\t/a/aludat [13],\t/a/aludat [13]}),
    .b({_al_u2697_o,_al_u2697_o}),
    .c({_al_u2614_o,_al_u2614_o}),
    .d({_al_u2616_o,_al_u2616_o}),
    .mi({open_n14371,\t/a/ID_read_dat1 [13]}),
    .fx({open_n14376,\t/a/ID_jump_regdat1 [13]}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2702|t/a/regfile/reg0_b1004  (
    .a({\t/a/aludat [12],_al_u2614_o}),
    .b({_al_u2701_o,_al_u2616_o}),
    .c({_al_u2614_o,\t/a/MEM_aludat [12]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [12]}),
    .e({\t/a/ID_read_dat1 [12],open_n14379}),
    .mi({open_n14381,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [12],_al_u2701_o}),
    .q({open_n14396,\t/a/regfile/regfile$31$ [12]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2706|t/a/regfile/reg0_b1003  (
    .a({\t/a/aludat [11],_al_u2614_o}),
    .b({_al_u2705_o,_al_u2616_o}),
    .c({_al_u2614_o,\t/a/MEM_aludat [11]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [11]}),
    .e({\t/a/ID_read_dat1 [11],open_n14397}),
    .mi({open_n14399,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [11],_al_u2705_o}),
    .q({open_n14414,\t/a/regfile/regfile$31$ [11]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~(~0*A))"),
    //.LUT1("(D*~C*~B*~(~1*A))"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000001100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2708 (
    .a({\t/a/alu/n5 [10],\t/a/alu/n5 [10]}),
    .b({_al_u2707_o,_al_u2707_o}),
    .c({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .d({_al_u2128_o,_al_u2128_o}),
    .mi({open_n14427,\t/a/EX_operation [0]}),
    .fx({open_n14432,_al_u2708_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(~0*~(~B*A))))"),
    //.LUTF1("~(~D*~(C*~(~0*~(~B*A))))"),
    //.LUTG0("~(~D*~(C*~(~1*~(~B*A))))"),
    //.LUTG1("~(~D*~(C*~(~1*~(~B*A))))"),
    .INIT_LUTF0(16'b1111111100100000),
    .INIT_LUTF1(16'b1111111100100000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2712|_al_u2715  (
    .a({_al_u2709_o,_al_u2709_o}),
    .b({_al_u2486_o,_al_u2486_o}),
    .c({_al_u2710_o,_al_u2713_o}),
    .d({_al_u2711_o,_al_u2714_o}),
    .e({_al_u2610_o,_al_u2616_o}),
    .f({\t/a/ID_jump_regdat2 [10],\t/a/ID_jump_regdat1 [10]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2717 (
    .a({\t/a/aludat [9],\t/a/aludat [9]}),
    .b({_al_u2716_o,_al_u2716_o}),
    .c({_al_u2606_o,_al_u2606_o}),
    .d({_al_u2610_o,_al_u2610_o}),
    .mi({open_n14469,\t/a/ID_read_dat2 [9]}),
    .fx({open_n14474,\t/a/ID_jump_regdat2 [9]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(0*~(D)*~(A)+0*D*~(A)+~(0)*D*A+0*D*A)))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(C*~(B*~(1*~(D)*~(A)+1*D*~(A)+~(1)*D*A+1*D*A)))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUTF0(16'b1011000000110000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1111000001110000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2719|_al_u1065  (
    .a({\t/a/aludat [9],\t/a/ID_rs2 [0]}),
    .b({_al_u2718_o,\t/a/ID_rs2 [1]}),
    .c({_al_u2614_o,\t/a/ID_rs2 [2]}),
    .d({_al_u2616_o,\t/a/regfile/regfile$31$ [9]}),
    .e({\t/a/ID_read_dat1 [9],\t/a/regfile/regfile$30$ [9]}),
    .f({\t/a/ID_jump_regdat1 [9],_al_u1065_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2721|t/a/regfile/reg0_b136  (
    .a({\t/a/aludat [8],_al_u2606_o}),
    .b({_al_u2720_o,_al_u2610_o}),
    .c({_al_u2606_o,\t/a/MEM_aludat [8]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o,\t/a/reg_writedat [8]}),
    .e({\t/a/ID_read_dat2 [8],open_n14499}),
    .mi({open_n14501,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [8],_al_u2720_o}),
    .q({open_n14516,\t/a/regfile/regfile$4$ [8]}));  // register.v(63)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2723|t/a/id_ex/reg8_b8  (
    .a({\t/a/aludat [8],_al_u333_o}),
    .b({_al_u2722_o,_al_u364_o}),
    .c({_al_u2614_o,_al_u374_o}),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [8]}),
    .e({\t/a/ID_read_dat1 [8],open_n14518}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [8],\t/a/ID_read_dat1 [8]}),
    .q({open_n14536,\t/a/EX_regdat1 [8]}));  // flow_line_reg.v(139)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2725|t/a/regfile/reg0_b135  (
    .a({\t/a/aludat [7],_al_u2606_o}),
    .b({_al_u2724_o,_al_u2610_o}),
    .c({_al_u2606_o,\t/a/MEM_aludat [7]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o,\t/a/reg_writedat [7]}),
    .e({\t/a/ID_read_dat2 [7],open_n14537}),
    .mi({open_n14539,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [7],_al_u2724_o}),
    .q({open_n14554,\t/a/regfile/regfile$4$ [7]}));  // register.v(63)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2727|t/a/id_ex/reg8_b7  (
    .a({\t/a/aludat [7],_al_u333_o}),
    .b({_al_u2726_o,_al_u385_o}),
    .c({_al_u2614_o,_al_u395_o}),
    .clk(clock_pad),
    .d({_al_u2616_o,\t/a/reg_writedat [7]}),
    .e({\t/a/ID_read_dat1 [7],open_n14556}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [7],\t/a/ID_read_dat1 [7]}),
    .q({open_n14574,\t/a/EX_regdat1 [7]}));  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUTF1("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUTG0("~(~D*~(C*~(~1*~(B*~A))))"),
    //.LUTG1("~(~D*~(C*~(~1*~(B*~A))))"),
    .INIT_LUTF0(16'b1111111101000000),
    .INIT_LUTF1(16'b1111111101000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111111111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2731|_al_u2734  (
    .a({_al_u2728_o,_al_u2728_o}),
    .b({_al_u2525_o,_al_u2525_o}),
    .c({_al_u2729_o,_al_u2732_o}),
    .d({_al_u2730_o,_al_u2733_o}),
    .e({_al_u2610_o,_al_u2616_o}),
    .f({\t/a/ID_jump_regdat2 [6],\t/a/ID_jump_regdat1 [6]}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2732|t/a/id_ex/reg8_b6  (
    .a({open_n14597,_al_u333_o}),
    .b({_al_u2616_o,_al_u406_o}),
    .c({\t/a/ID_read_dat1 [6],_al_u416_o}),
    .clk(clock_pad),
    .d({_al_u2614_o,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u2732_o,\t/a/ID_read_dat1 [6]}),
    .q({open_n14614,\t/a/EX_regdat1 [6]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(~(A)*~(B)*~(D)+~(A)*~(B)*D+A*~(B)*D+~(A)*B*D))"),
    //.LUT1("(D*~(~B*~(~C*~A)))"),
    .INIT_LUT0(16'b0111000000010000),
    .INIT_LUT1(16'b1100110100000000),
    .MODE("LOGIC"))
    \_al_u2735|_al_u2536  (
    .a({\t/a/alu/mux0_b5/B1_0 ,\t/a/EX_A [5]}),
    .b({_al_u2536_o,\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o }),
    .c(\t/a/EX_operation [2:1]),
    .d({_al_u2128_o,\t/a/EX_operation [0]}),
    .f({_al_u2735_o,_al_u2536_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("~(~D*~(C*~(~1*~(B*~A))))"),
    //.LUTG1("(D*~(~C*B))"),
    .INIT_LUTF0(16'b1111111101000000),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2736|_al_u2738  (
    .a({open_n14635,_al_u2735_o}),
    .b({_al_u2610_o,_al_u2535_o}),
    .c({\t/a/ID_read_dat2 [5],_al_u2736_o}),
    .d({_al_u2606_o,_al_u2737_o}),
    .e({open_n14638,_al_u2610_o}),
    .f({_al_u2736_o,\t/a/ID_jump_regdat2 [5]}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2739|t/a/id_ex/reg8_b5  (
    .a({open_n14659,_al_u333_o}),
    .b({_al_u2616_o,_al_u427_o}),
    .c({\t/a/ID_read_dat1 [5],_al_u437_o}),
    .clk(clock_pad),
    .d({_al_u2614_o,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u2739_o,\t/a/ID_read_dat1 [5]}),
    .q({open_n14676,\t/a/EX_regdat1 [5]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(B*~A))))"),
    .INIT_LUT0(16'b1111111101000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2741 (
    .a({_al_u2735_o,_al_u2735_o}),
    .b({_al_u2535_o,_al_u2535_o}),
    .c({_al_u2739_o,_al_u2739_o}),
    .d({_al_u2740_o,_al_u2740_o}),
    .mi({open_n14689,_al_u2616_o}),
    .fx({open_n14694,\t/a/ID_jump_regdat1 [5]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2743 (
    .a({\t/a/aludat [4],\t/a/aludat [4]}),
    .b({_al_u2742_o,_al_u2742_o}),
    .c({_al_u2606_o,_al_u2606_o}),
    .d({_al_u2610_o,_al_u2610_o}),
    .mi({open_n14709,\t/a/ID_read_dat2 [4]}),
    .fx({open_n14714,\t/a/ID_jump_regdat2 [4]}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTF1("(D*~(~C*B))"),
    //.LUTG0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG1("(D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101100000001),
    .INIT_LUTF1(16'b1111001100000000),
    .INIT_LUTG0(16'b1010101100000001),
    .INIT_LUTG1(16'b1111001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2744|t/a/id_ex/reg8_b4  (
    .a({open_n14717,_al_u333_o}),
    .b({_al_u2616_o,_al_u448_o}),
    .c({\t/a/ID_read_dat1 [4],_al_u458_o}),
    .clk(clock_pad),
    .d({_al_u2614_o,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u2744_o,\t/a/ID_read_dat1 [4]}),
    .q({open_n14738,\t/a/EX_regdat1 [4]}));  // flow_line_reg.v(139)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("~(~B*~((~D*~C))*~(A)+~B*(~D*~C)*~(A)+~(~B)*(~D*~C)*A+~B*(~D*~C)*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b1110111011100100),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2746|t/a/regfile/reg0_b132  (
    .a({_al_u2744_o,_al_u2614_o}),
    .b({_al_u2745_o,_al_u2616_o}),
    .c({_al_u2616_o,\t/a/MEM_aludat [4]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/aludat [4],\t/a/reg_writedat [4]}),
    .mi({open_n14749,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat1 [4],_al_u2745_o}),
    .q({open_n14753,\t/a/regfile/regfile$4$ [4]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*(~(A)*~(B)*~(D)+~(A)*~(B)*D+A*~(B)*D+~(A)*B*D))"),
    //.LUT1("(D*~(~B*~(~C*~A)))"),
    .INIT_LUT0(16'b0111000000010000),
    .INIT_LUT1(16'b1100110100000000),
    .MODE("LOGIC"))
    \_al_u2747|_al_u2556  (
    .a({\t/a/alu/mux0_b3/B1_0 ,\t/a/EX_A [3]}),
    .b({_al_u2556_o,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .c(\t/a/EX_operation [2:1]),
    .d({_al_u2128_o,\t/a/EX_operation [0]}),
    .f({_al_u2747_o,_al_u2556_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(B*~A))))"),
    .INIT_LUT0(16'b1111111101000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2750 (
    .a({_al_u2747_o,_al_u2747_o}),
    .b({_al_u2555_o,_al_u2555_o}),
    .c({_al_u2748_o,_al_u2748_o}),
    .d({_al_u2749_o,_al_u2749_o}),
    .mi({open_n14786,_al_u2610_o}),
    .fx({open_n14791,\t/a/ID_jump_regdat2 [3]}));
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("(D*~(~C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1111001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2751|t/a/id_ex/reg8_b3  (
    .a({open_n14794,_al_u333_o}),
    .b({_al_u2616_o,_al_u469_o}),
    .c({\t/a/ID_read_dat1 [3],_al_u479_o}),
    .clk(clock_pad),
    .d({_al_u2614_o,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u2751_o,\t/a/ID_read_dat1 [3]}),
    .q({open_n14811,\t/a/EX_regdat1 [3]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(B*~A))))"),
    .INIT_LUT0(16'b1111111101000000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2753 (
    .a({_al_u2747_o,_al_u2747_o}),
    .b({_al_u2555_o,_al_u2555_o}),
    .c({_al_u2751_o,_al_u2751_o}),
    .d({_al_u2752_o,_al_u2752_o}),
    .mi({open_n14824,_al_u2616_o}),
    .fx({open_n14829,\t/a/ID_jump_regdat1 [3]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2755|_al_u2757  (
    .a({\t/a/aludat [2],\t/a/aludat [2]}),
    .b({_al_u2754_o,_al_u2756_o}),
    .c({_al_u2606_o,_al_u2614_o}),
    .d({_al_u2610_o,_al_u2616_o}),
    .e({\t/a/ID_read_dat2 [2],\t/a/ID_read_dat1 [2]}),
    .f({\t/a/ID_jump_regdat2 [2],\t/a/ID_jump_regdat1 [2]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2759|_al_u2761  (
    .a({\t/a/aludat [0],\t/a/aludat [0]}),
    .b({_al_u2758_o,_al_u2760_o}),
    .c({_al_u2606_o,_al_u2614_o}),
    .d({_al_u2610_o,_al_u2616_o}),
    .e({\t/a/ID_read_dat2 [0],\t/a/ID_read_dat1 [0]}),
    .f({\t/a/ID_jump_regdat2 [0],\t/a/ID_jump_regdat1 [0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*~A)"),
    //.LUT1("(~1*~D*~C*~B*~A)"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u276 (
    .a({\t/a/WB_rd [0],\t/a/WB_rd [0]}),
    .b({\t/a/WB_rd [1],\t/a/WB_rd [1]}),
    .c({\t/a/WB_rd [2],\t/a/WB_rd [2]}),
    .d({\t/a/WB_rd [3],\t/a/WB_rd [3]}),
    .mi({open_n14888,\t/a/WB_rd [4]}),
    .fx({open_n14893,\t/a/regfile/n46 [0]}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTF1("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTG0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000101000000),
    .INIT_LUTF1(16'b1100110011101100),
    .INIT_LUTG0(16'b0101000101000000),
    .INIT_LUTG1(16'b1111110011101100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2763|t/a/regfile/reg0_b129  (
    .a({\t/a/aludat [1],_al_u2606_o}),
    .b({_al_u2762_o,_al_u2610_o}),
    .c({_al_u2606_o,\t/a/MEM_aludat [1]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({_al_u2610_o,\t/a/reg_writedat [1]}),
    .e({\t/a/ID_read_dat2 [1],open_n14896}),
    .mi({open_n14898,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({\t/a/ID_jump_regdat2 [1],_al_u2762_o}),
    .q({open_n14913,\t/a/regfile/regfile$4$ [1]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUT1("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    .INIT_LUT0(16'b1100110011101100),
    .INIT_LUT1(16'b1111110011101100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2765 (
    .a({\t/a/aludat [1],\t/a/aludat [1]}),
    .b({_al_u2764_o,_al_u2764_o}),
    .c({_al_u2614_o,_al_u2614_o}),
    .d({_al_u2616_o,_al_u2616_o}),
    .mi({open_n14926,\t/a/ID_read_dat1 [1]}),
    .fx({open_n14931,\t/a/ID_jump_regdat1 [1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~C)*~(B@A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(D*~C)*~(B@A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1001000010011001),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1001000010011001),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2767|_al_u2770  (
    .a({open_n14934,\t/a/ID_jump_regdat2 [14]}),
    .b({open_n14935,\t/a/ID_jump_regdat1 [14]}),
    .c({\t/a/ID_jump_regdat1 [1],\t/a/ID_jump_regdat2 [1]}),
    .d({\t/a/ID_jump_regdat2 [1],\t/a/ID_jump_regdat1 [1]}),
    .f({_al_u2767_o,_al_u2770_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0@D)*~(C@B))"),
    //.LUT1("(~A*~(1@D)*~(C@B))"),
    .INIT_LUT0(16'b0000000001000001),
    .INIT_LUT1(16'b0100000100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2768 (
    .a({_al_u2767_o,_al_u2767_o}),
    .b({\t/a/ID_jump_regdat2 [13],\t/a/ID_jump_regdat2 [13]}),
    .c({\t/a/ID_jump_regdat1 [13],\t/a/ID_jump_regdat1 [13]}),
    .d({\t/a/ID_jump_regdat2 [4],\t/a/ID_jump_regdat2 [4]}),
    .mi({open_n14972,\t/a/ID_jump_regdat1 [4]}),
    .fx({open_n14977,_al_u2768_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("(~(D@C)*~(B@A))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("(~(D@C)*~(B@A))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1001000000001001),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1001000000001001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2769|_al_u2668  (
    .a({\t/a/ID_jump_regdat2 [18],\t/a/aludat [18]}),
    .b({\t/a/ID_jump_regdat1 [18],_al_u2667_o}),
    .c({\t/a/ID_jump_regdat2 [5],_al_u2606_o}),
    .d({\t/a/ID_jump_regdat1 [5],_al_u2610_o}),
    .e({open_n14982,\t/a/ID_read_dat2 [18]}),
    .f({_al_u2769_o,\t/a/ID_jump_regdat2 [18]}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D*~C)*~(B*~A))"),
    //.LUT1("(~(D@C)*~(B@A))"),
    .INIT_LUT0(16'b1011000010111011),
    .INIT_LUT1(16'b1001000000001001),
    .MODE("LOGIC"))
    \_al_u2772|_al_u2776  (
    .a({\t/a/ID_jump_regdat2 [22],\t/a/ID_jump_regdat2 [28]}),
    .b({\t/a/ID_jump_regdat1 [22],\t/a/ID_jump_regdat1 [28]}),
    .c({\t/a/ID_jump_regdat2 [21],\t/a/ID_jump_regdat2 [26]}),
    .d({\t/a/ID_jump_regdat1 [21],\t/a/ID_jump_regdat1 [26]}),
    .f({_al_u2772_o,_al_u2776_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(B*A*~(D@C))"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2773|_al_u2771  (
    .a({_al_u2771_o,_al_u2768_o}),
    .b({_al_u2772_o,_al_u2769_o}),
    .c({\t/a/ID_jump_regdat2 [31],_al_u2770_o}),
    .d({\t/a/ID_jump_regdat1 [31],\t/a/ID_jump_regdat2 [10]}),
    .e({open_n15025,\t/a/ID_jump_regdat1 [10]}),
    .f({_al_u2773_o,_al_u2771_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2774|_al_u2636  (
    .a({open_n15046,\t/a/aludat [26]}),
    .b({open_n15047,_al_u2635_o}),
    .c({\t/a/ID_jump_regdat1 [26],_al_u2606_o}),
    .d({\t/a/ID_jump_regdat2 [26],_al_u2610_o}),
    .e({open_n15050,\t/a/ID_read_dat2 [26]}),
    .f({_al_u2774_o,\t/a/ID_jump_regdat2 [26]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@D)*~(~C*B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(~A*~(1@D)*~(~C*B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .INIT_LUTF0(16'b0000000001010001),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0101000100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2777|_al_u2775  (
    .a({_al_u2773_o,_al_u2774_o}),
    .b({_al_u2775_o,\t/a/ID_jump_regdat2 [28]}),
    .c({_al_u2776_o,\t/a/ID_jump_regdat1 [28]}),
    .d({\t/a/ID_jump_regdat2 [19],\t/a/ID_jump_regdat2 [24]}),
    .e({\t/a/ID_jump_regdat1 [19],\t/a/ID_jump_regdat1 [24]}),
    .f({_al_u2777_o,_al_u2775_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("(~(D@C)*~(B@A))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("(~(D@C)*~(B@A))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1001000000001001),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1001000000001001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2778|_al_u2620  (
    .a({\t/a/ID_jump_regdat2 [30],\t/a/aludat [30]}),
    .b({\t/a/ID_jump_regdat1 [30],_al_u2619_o}),
    .c({\t/a/ID_jump_regdat2 [25],_al_u2606_o}),
    .d({\t/a/ID_jump_regdat1 [25],_al_u2610_o}),
    .e({open_n15095,\t/a/ID_read_dat2 [30]}),
    .f({_al_u2778_o,\t/a/ID_jump_regdat2 [30]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("(A*~(0@D)*~(C@B))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("(A*~(1@D)*~(C@B))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b0000000010000010),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1000001000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2779|_al_u2624  (
    .a({_al_u2778_o,\t/a/aludat [29]}),
    .b({\t/a/ID_jump_regdat2 [29],_al_u2623_o}),
    .c({\t/a/ID_jump_regdat1 [29],_al_u2606_o}),
    .d({\t/a/ID_jump_regdat2 [27],_al_u2610_o}),
    .e({\t/a/ID_jump_regdat1 [27],\t/a/ID_read_dat2 [29]}),
    .f({_al_u2779_o,\t/a/ID_jump_regdat2 [29]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D@C)*~(B*~A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(D@C)*~(B*~A))"),
    //.LUTG1("(~C*D)"),
    .INIT_LUTF0(16'b1011000000001011),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1011000000001011),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2780|_al_u2782  (
    .a({open_n15138,\t/a/ID_jump_regdat2 [6]}),
    .b({open_n15139,\t/a/ID_jump_regdat1 [6]}),
    .c({\t/a/ID_jump_regdat1 [6],\t/a/ID_jump_regdat2 [2]}),
    .d({\t/a/ID_jump_regdat2 [6],\t/a/ID_jump_regdat1 [2]}),
    .f({_al_u2780_o,_al_u2782_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("(~A*~(0@D)*~(C*~B))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("(~A*~(1@D)*~(C*~B))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b0000000001000101),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b0100010100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2781|_al_u2672  (
    .a({_al_u2780_o,\t/a/aludat [17]}),
    .b({\t/a/ID_jump_regdat2 [20],_al_u2671_o}),
    .c({\t/a/ID_jump_regdat1 [20],_al_u2606_o}),
    .d({\t/a/ID_jump_regdat2 [17],_al_u2610_o}),
    .e({\t/a/ID_jump_regdat1 [17],\t/a/ID_read_dat2 [17]}),
    .f({_al_u2781_o,\t/a/ID_jump_regdat2 [17]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("(B*A*~(D@C))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2783|_al_u2650  (
    .a({_al_u2781_o,\t/a/aludat [23]}),
    .b({_al_u2782_o,_al_u2649_o}),
    .c({\t/a/ID_jump_regdat2 [23],_al_u2614_o}),
    .d({\t/a/ID_jump_regdat1 [23],_al_u2616_o}),
    .e({open_n15188,\t/a/ID_read_dat1 [23]}),
    .f({_al_u2783_o,\t/a/ID_jump_regdat1 [23]}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("(~(D@C)*~(B@A))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("(~(D@C)*~(B@A))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b1001000000001001),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b1001000000001001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2784|_al_u2700  (
    .a({\t/a/ID_jump_regdat2 [12],\t/a/aludat [12]}),
    .b({\t/a/ID_jump_regdat1 [12],_al_u2699_o}),
    .c({\t/a/ID_jump_regdat2 [8],_al_u2606_o}),
    .d({\t/a/ID_jump_regdat1 [8],_al_u2610_o}),
    .e({open_n15211,\t/a/ID_read_dat2 [12]}),
    .f({_al_u2784_o,\t/a/ID_jump_regdat2 [12]}));
  EG_PHY_MSLICE #(
    //.LUT0("(A*~(0@D)*~(C@B))"),
    //.LUT1("(A*~(1@D)*~(C@B))"),
    .INIT_LUT0(16'b0000000010000010),
    .INIT_LUT1(16'b1000001000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2787 (
    .a({_al_u2786_o,_al_u2786_o}),
    .b({\t/a/ID_jump_regdat2 [0],\t/a/ID_jump_regdat2 [0]}),
    .c({\t/a/ID_jump_regdat1 [0],\t/a/ID_jump_regdat1 [0]}),
    .d({\t/a/ID_jump_regdat2 [9],\t/a/ID_jump_regdat2 [9]}),
    .mi({open_n15244,\t/a/ID_jump_regdat1 [9]}),
    .fx({open_n15249,_al_u2787_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~(D@C)*~(~B*A))"),
    //.LUT1("(C*~D)"),
    .INIT_LUT0(16'b1101000000001101),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"))
    \_al_u2788|_al_u2786  (
    .a({open_n15252,\t/a/ID_jump_regdat2 [15]}),
    .b({open_n15253,\t/a/ID_jump_regdat1 [15]}),
    .c({\t/a/ID_jump_regdat1 [15],\t/a/ID_jump_regdat2 [7]}),
    .d({\t/a/ID_jump_regdat2 [15],\t/a/ID_jump_regdat1 [7]}),
    .f({_al_u2788_o,_al_u2786_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~(~B*~(C*(A*~(0)*~(D)+A*0*~(D)+~(A)*0*D+A*0*D)))"),
    //.LUTF1("(~A*~(0@D)*~(C@B))"),
    //.LUTG0("~(~B*~(C*(A*~(1)*~(D)+A*1*~(D)+~(A)*1*D+A*1*D)))"),
    //.LUTG1("(~A*~(1@D)*~(C@B))"),
    .INIT_LUTF0(16'b1100110011101100),
    .INIT_LUTF1(16'b0000000001000001),
    .INIT_LUTG0(16'b1111110011101100),
    .INIT_LUTG1(16'b0100000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2789|_al_u2704  (
    .a({_al_u2788_o,\t/a/aludat [11]}),
    .b({\t/a/ID_jump_regdat2 [11],_al_u2703_o}),
    .c({\t/a/ID_jump_regdat1 [11],_al_u2606_o}),
    .d({\t/a/ID_jump_regdat2 [3],_al_u2610_o}),
    .e({\t/a/ID_jump_regdat1 [3],\t/a/ID_read_dat2 [11]}),
    .f({_al_u2789_o,\t/a/ID_jump_regdat2 [11]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(0@D)*~(~C*B))"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(A*~(1@D)*~(~C*B))"),
    //.LUTG1("(1*D*C*B*A)"),
    .INIT_LUTF0(16'b0000000010100010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010001000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2790|_al_u2785  (
    .a({_al_u2779_o,_al_u2784_o}),
    .b({_al_u2783_o,\t/a/ID_jump_regdat2 [20]}),
    .c({_al_u2785_o,\t/a/ID_jump_regdat1 [20]}),
    .d({_al_u2787_o,\t/a/ID_jump_regdat2 [16]}),
    .e({_al_u2789_o,\t/a/ID_jump_regdat1 [16]}),
    .f({_al_u2790_o,_al_u2785_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("(~D*~(C*~(~B*~A)))"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("(~D*~(C*~(~B*~A)))"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0000000000011111),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0000000000011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2792|_al_u1756  (
    .a({_al_u2766_o,\t/a/condition/n5 [4]}),
    .b({_al_u2791_o,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/n1_lutinv ,\t/a/condition/n1_lutinv }),
    .d({\t/a/condition/sel1/B2 ,\t/a/condition/sel1/B2 }),
    .e({open_n15320,\t/a/ID_rd [4]}),
    .f({_al_u2792_o,\t/a/ID_jump_addr [4]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("(~(~C*~B)*~(D*A))"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("(~(~C*~B)*~(D*A))"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0101010011111100),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0101010011111100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2794|_al_u1782  (
    .a({_al_u1958_o,\t/a/condition/n5 [1]}),
    .b({_al_u1965_o,\t/a/condition/n0_lutinv }),
    .c({\t/a/ID_rd [1],\t/a/condition/n1_lutinv }),
    .d({\t/a/ID_rd [3],\t/a/condition/sel1/B2 }),
    .e({open_n15343,\t/a/ID_rd [1]}),
    .f({_al_u2794_o,\t/a/ID_jump_addr [1]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("(~(C*B)*~(~D*~A))"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("(~(C*B)*~(~D*~A))"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0011111100101010),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0011111100101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2795|_al_u1760  (
    .a({_al_u1958_o,\t/a/condition/n5 [3]}),
    .b({_al_u1962_o,\t/a/condition/n0_lutinv }),
    .c({\t/a/ID_rd [0],\t/a/condition/n1_lutinv }),
    .d({\t/a/ID_rd [3],\t/a/condition/sel1/B2 }),
    .e({open_n15366,\t/a/ID_rd [3]}),
    .f({_al_u2795_o,\t/a/ID_jump_addr [3]}));
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(~C*B))"),
    //.LUT1("(~(D*B)*~(~C*~A))"),
    .INIT_LUT0(16'b1111111100001100),
    .INIT_LUT1(16'b0011001011111010),
    .MODE("LOGIC"))
    \_al_u2796|_al_u2091  (
    .a({_al_u1962_o,open_n15387}),
    .b({_al_u1965_o,_al_u2080_o}),
    .c({\t/a/ID_rd [0],_al_u1962_o}),
    .d({\t/a/ID_rd [1],_al_u2078_o}),
    .f({_al_u2796_o,\t/a/IF_skip_addr [20]}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(D*C*B*A)"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2797|_al_u1742  (
    .a({_al_u2793_o,open_n15408}),
    .b({_al_u2794_o,open_n15409}),
    .c({_al_u2795_o,\t/a/ID_rs1 [2]}),
    .d({_al_u2796_o,\t/a/EX_rd [2]}),
    .f({\t/a/n4_lutinv ,_al_u1742_o}));
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(~C*~B)*~(~D*~A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(~C*~B)*~(~D*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1111110010101000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1111110010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2798|t/a/id_ex/reg5_b1  (
    .a({_al_u2113_o,open_n15434}),
    .b({_al_u2117_o,open_n15435}),
    .c({\t/a/ID_rd [1],\t/a/ID_rd [1]}),
    .clk(clock_pad),
    .d({\t/a/ID_rd [3],_al_u2117_o}),
    .mi({open_n15440,\t/a/ID_rd [1]}),
    .sr(rst_pad),
    .f({_al_u2798_o,_al_u2800_o}),
    .q({open_n15455,\t/a/EX_rd [1]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2802|t/a/if_id/reg6_b3  (
    .c({\t/instruction$3$_neg_lutinv ,\t/instruction$3$_neg_lutinv }),
    .clk(clock_pad),
    .d({\t/instruction$2$_neg_lutinv ,\t/a/if_id/n9 }),
    .sr(rst_pad),
    .f({_al_u2802_o,open_n15473}),
    .q({open_n15477,\t/a/ID_op [3]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~B*A*(0@D))"),
    //.LUTF1("(0*~(C*~(~A*~(D*B))))"),
    //.LUTG0("(~C*~B*A*(1@D))"),
    //.LUTG1("(1*~(C*~(~A*~(D*B))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b0001111101011111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2807|t/a/id_ex/reg5_b2  (
    .a({\t/a/n4_lutinv ,_al_u2798_o}),
    .b({_al_u2801_o,_al_u2799_o}),
    .c({\t/a/n2 ,_al_u2800_o}),
    .clk(clock_pad),
    .d({_al_u2806_o,_al_u2115_o}),
    .e({\t/busarbitration/n3 ,\t/a/ID_rd [2]}),
    .mi({open_n15480,\t/a/ID_rd [2]}),
    .sr(rst_pad),
    .f({_al_u2807_o,_al_u2801_o}),
    .q({open_n15495,\t/a/EX_rd [2]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111100010),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1111001111100010),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2808|t/a/id_ex/reg7_b9  (
    .a({open_n15496,_al_u2807_o}),
    .b({open_n15497,\t/a/condition/n0_lutinv }),
    .c({\t/a/condition/n0_lutinv ,\t/a/ID_memstraddr [9]}),
    .clk(clock_pad),
    .d({_al_u2807_o,\t/memstraddress [9]}),
    .mi({open_n15502,\t/a/ID_memstraddr [9]}),
    .sr(rst_pad),
    .f({_al_u2808_o,_al_u2812_o}),
    .q({open_n15517,\t/a/EX_memstraddr [9]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("~(~C*B*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("~(~C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111001111111111),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111001111111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u2809|t/a/if_id/reg5_b18  (
    .b({_al_u2808_o,\t/a/MEM_aludat [18]}),
    .c({\t/instrnop ,\t/memstraddress [18]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({_al_u2792_o,\t/busarbitration/n3 }),
    .mi({open_n15523,\t/memstraddress [18]}),
    .sr(rst_pad),
    .f({\t/a/if_id/n9 ,addr[18]}),
    .q({open_n15538,\t/a/ID_memstraddr [18]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b1011000010000000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1011000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2811|_al_u2880  (
    .a({n8[8],n8[11]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,\t/a/instr/n12 [12]}),
    .d({\t/a/instr/n16 [7],_al_u2109_o}),
    .e({open_n15541,\t/a/instr/n16 [10]}),
    .f({_al_u2811_o,_al_u2880_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b1011000010000000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1011000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2814|_al_u2866  (
    .a({n8[7],n8[16]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,\t/a/instr/n12 [17]}),
    .d({\t/a/instr/n16 [6],_al_u2109_o}),
    .e({open_n15564,\t/a/instr/n16 [15]}),
    .f({_al_u2814_o,_al_u2866_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b1000100011110000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1011101111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2817|_al_u2854  (
    .a({n8[6],n8[20]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [7],\t/a/instr/n12 [21]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .e({\t/a/instr/n16 [5],\t/a/instr/n16 [19]}),
    .f({_al_u2817_o,_al_u2854_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b1000100011110000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1011101111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2819|_al_u2852  (
    .a({n8[5],n8[21]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [6],\t/a/instr/n12 [22]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .e({\t/a/instr/n16 [4],\t/a/instr/n16 [20]}),
    .f({_al_u2819_o,_al_u2852_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b1011000010000000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1011000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2821|_al_u2831  (
    .a({n8[4],n8[2]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,\t/a/instr/n12 [3]}),
    .d({\t/a/instr/n16 [3],_al_u2109_o}),
    .e({open_n15631,\t/a/instr/n16 [1]}),
    .f({_al_u2821_o,_al_u2831_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTF1("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUTG0("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    //.LUTG1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUTF0(16'b1000100011110000),
    .INIT_LUTF1(16'b1000100011110000),
    .INIT_LUTG0(16'b1011101111110000),
    .INIT_LUTG1(16'b1011101111110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2824|_al_u2826  (
    .a({n8[3],n8[30]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [4],\t/a/instr/n12 [31]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .e({\t/a/instr/n16 [2],\t/a/instr/n16 [29]}),
    .f({_al_u2824_o,_al_u2826_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1011000010000000),
    .MODE("LOGIC"))
    \_al_u2828|_al_u2110  (
    .a({n8[29],_al_u2109_o}),
    .b({_al_u2810_o,\t/busarbitration/n3 }),
    .c({_al_u2109_o,\t/busarbitration/instruction [31]}),
    .d({\t/a/instr/n16 [28],i_data[31]}),
    .f({_al_u2828_o,\t/a/IF_skip_addr [31]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    //.LUT1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUT0(16'b1101000010000000),
    .INIT_LUT1(16'b1011000010000000),
    .MODE("LOGIC"))
    \_al_u2833|_al_u2887  (
    .a({n8[28],_al_u2810_o}),
    .b({_al_u2810_o,n8[0]}),
    .c({_al_u2109_o,_al_u2109_o}),
    .d({\t/a/instr/n16 [27],\t/memstraddress [1]}),
    .f({_al_u2833_o,_al_u2887_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUT1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUT0(16'b1000100011110000),
    .INIT_LUT1(16'b1011101111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2836 (
    .a({n8[27],n8[27]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [28],\t/a/instr/n12 [28]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .mi({open_n15726,\t/a/instr/n16 [26]}),
    .fx({open_n15731,_al_u2836_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUT1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUT0(16'b1000100011110000),
    .INIT_LUT1(16'b1011101111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2838 (
    .a({n8[26],n8[26]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [27],\t/a/instr/n12 [27]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .mi({open_n15746,\t/a/instr/n16 [25]}),
    .fx({open_n15751,_al_u2838_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~D)"),
    //.LUT1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUT0(16'b0000000000001111),
    .INIT_LUT1(16'b1011000010000000),
    .MODE("LOGIC"))
    \_al_u2840|_al_u2810  (
    .a({n8[25],open_n15754}),
    .b({_al_u2810_o,open_n15755}),
    .c({_al_u2109_o,\t/a/condition/n0_lutinv }),
    .d({\t/a/instr/n16 [24],_al_u2792_o}),
    .f({_al_u2840_o,_al_u2810_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTF1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTG0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTG1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUTF0(16'b1011000010000000),
    .INIT_LUTF1(16'b1011000010000000),
    .INIT_LUTG0(16'b1011000010000000),
    .INIT_LUTG1(16'b1011000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2843|_al_u2882  (
    .a({n8[24],n8[10]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,_al_u2109_o}),
    .d({\t/a/instr/n16 [23],\t/a/instr/n16 [9]}),
    .f({_al_u2843_o,_al_u2882_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTF1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTG0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTG1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUTF0(16'b1011000010000000),
    .INIT_LUTF1(16'b1011000010000000),
    .INIT_LUTG0(16'b1011000010000000),
    .INIT_LUTG1(16'b1011000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2846|_al_u2877  (
    .a({n8[23],n8[12]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,_al_u2109_o}),
    .d({\t/a/instr/n16 [22],\t/a/instr/n16 [11]}),
    .f({_al_u2846_o,_al_u2877_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUT1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUT0(16'b1011000010000000),
    .INIT_LUT1(16'b1011000010000000),
    .MODE("LOGIC"))
    \_al_u2849|_al_u2874  (
    .a({n8[22],n8[13]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,_al_u2109_o}),
    .d({\t/a/instr/n16 [21],\t/a/instr/n16 [12]}),
    .f({_al_u2849_o,_al_u2874_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUT1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUT0(16'b1011000010000000),
    .INIT_LUT1(16'b1011000010000000),
    .MODE("LOGIC"))
    \_al_u2856|_al_u2871  (
    .a({n8[19],n8[14]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,_al_u2109_o}),
    .d({\t/a/instr/n16 [18],\t/a/instr/n16 [13]}),
    .f({_al_u2856_o,_al_u2871_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTF1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTG0("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    //.LUTG1("(C*(D*~(A)*~(B)+D*A*~(B)+~(D)*A*B+D*A*B))"),
    .INIT_LUTF0(16'b1011000010000000),
    .INIT_LUTF1(16'b1011000010000000),
    .INIT_LUTG0(16'b1011000010000000),
    .INIT_LUTG1(16'b1011000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2859|_al_u2868  (
    .a({n8[1],n8[15]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({_al_u2109_o,_al_u2109_o}),
    .d({\t/a/instr/n16 [0],\t/a/instr/n16 [14]}),
    .f({_al_u2859_o,_al_u2868_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUT1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUT0(16'b1000100011110000),
    .INIT_LUT1(16'b1011101111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2862 (
    .a({n8[18],n8[18]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [19],\t/a/instr/n12 [19]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .mi({open_n15900,\t/a/instr/n16 [17]}),
    .fx({open_n15905,_al_u2862_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUT1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUT0(16'b1000100011110000),
    .INIT_LUT1(16'b1011101111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2864 (
    .a({n8[17],n8[17]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [18],\t/a/instr/n12 [18]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .mi({open_n15920,\t/a/instr/n16 [16]}),
    .fx({open_n15925,_al_u2864_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*~(D)+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)+~(C)*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D+C*(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D)"),
    //.LUT1("(C*~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*~(D)+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)+~(C)*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D+C*(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D)"),
    .INIT_LUT0(16'b1000100011110000),
    .INIT_LUT1(16'b1011101111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2885 (
    .a({n8[9],n8[9]}),
    .b({_al_u2810_o,_al_u2810_o}),
    .c({\t/a/instr/n12 [10],\t/a/instr/n12 [10]}),
    .d({_al_u2109_o,_al_u2109_o}),
    .mi({open_n15940,\t/a/instr/n16 [8]}),
    .fx({open_n15945,_al_u2885_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"))
    \_al_u322|_al_u1472  (
    .a({open_n15948,\t/a/ID_rs2 [0]}),
    .b({\t/a/MEM_aludat [1],\t/a/ID_rs2 [1]}),
    .c({\t/memstraddress [1],\t/a/regfile/regfile$0$ [1]}),
    .d({\t/busarbitration/n3 ,\t/a/regfile/regfile$1$ [1]}),
    .f({addr[1],_al_u1472_o}));
  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~((D*~B))*~(A)+C*(D*~B)*~(A)+~(C)*(D*~B)*A+C*(D*~B)*A)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111001001010000),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u323|t/a/mem_wb/reg0_b0  (
    .a({open_n15969,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .b({\t/a/MEM_aludat [0],_al_u1908_o}),
    .c({\t/memstraddress [0],\t/a/MEM_aludat [0]}),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,i_data[0]}),
    .sr(rst_pad),
    .f({addr[0],open_n15983}),
    .q({open_n15987,\t/a/reg_writedat [0]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u324|_al_u327  (
    .b({addr[5],addr[2]}),
    .c({memwrite_cs,memwrite_cs}),
    .d({n0,n0}),
    .f({n2[3],n2[0]}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"))
    \_al_u325|_al_u326  (
    .b(addr[4:3]),
    .c({memwrite_cs,memwrite_cs}),
    .d({n0,n0}),
    .f(n2[2:1]));
  EG_PHY_MSLICE #(
    //.LUT0("(~A*~(0@C)*~(D*~B))"),
    //.LUT1("(~A*~(1@C)*~(D*~B))"),
    .INIT_LUT0(16'b0000010000000101),
    .INIT_LUT1(16'b0100000001010000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u329 (
    .a({_al_u328_o,_al_u328_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [3],\t/a/ID_rs1 [3]}),
    .d({\t/a/WB_rd [0],\t/a/WB_rd [0]}),
    .mi({open_n16044,\t/a/WB_rd [3]}),
    .fx({open_n16049,_al_u329_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u330|_al_u359  (
    .a({\t/a/ID_rs1 [0],_al_u355_o}),
    .b({\t/a/ID_rs1 [4],_al_u356_o}),
    .c({\t/a/WB_rd [0],_al_u357_o}),
    .d({\t/a/WB_rd [4],_al_u358_o}),
    .e({open_n16054,\t/a/ID_rs1 [2]}),
    .f({_al_u330_o,_al_u359_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u331|_al_u915  (
    .a({\t/a/ID_rs1 [1],_al_u911_o}),
    .b({\t/a/ID_rs1 [4],_al_u912_o}),
    .c({\t/a/WB_rd [1],_al_u913_o}),
    .d({\t/a/WB_rd [4],_al_u914_o}),
    .e({open_n16077,\t/a/ID_rs1 [2]}),
    .f({_al_u331_o,_al_u915_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(C*B*A*~(0@D))"),
    //.LUT1("(C*B*A*~(1@D))"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u332 (
    .a({_al_u329_o,_al_u329_o}),
    .b({_al_u330_o,_al_u330_o}),
    .c({_al_u331_o,_al_u331_o}),
    .d({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .mi({open_n16110,\t/a/WB_rd [2]}),
    .fx({open_n16115,\t/a/regfile/n1_lutinv }));
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*~B*A)"),
    //.LUTF1("(C*D)"),
    //.LUTG0("(1*D*~C*~B*A)"),
    //.LUTG1("(C*D)"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1111000000000000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b1111000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u333|_al_u2613  (
    .a({open_n16118,\t/a/regfile/n1_lutinv }),
    .b({open_n16119,\t/a/risk_jump/n24_lutinv }),
    .c({\t/a/WB_regwritecs ,\t/a/risk_jump/n11_lutinv }),
    .d({\t/a/regfile/n1_lutinv ,\t/a/n19 }),
    .e({open_n16122,\t/a/condition/n1_lutinv }),
    .f({_al_u333_o,_al_u2613_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u338 (
    .a({_al_u334_o,_al_u334_o}),
    .b({_al_u335_o,_al_u335_o}),
    .c({_al_u336_o,_al_u336_o}),
    .d({_al_u337_o,_al_u337_o}),
    .mi({open_n16155,\t/a/ID_rs1 [2]}),
    .fx({open_n16160,_al_u338_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u343|t/a/regfile/reg0_b649  (
    .a({_al_u338_o,_al_u339_o}),
    .b({_al_u340_o,\t/a/ID_rs1 [0]}),
    .c({_al_u342_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [9]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [9]}),
    .mi({open_n16164,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u343_o,_al_u340_o}),
    .q({open_n16179,\t/a/regfile/regfile$20$ [9]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u344|_al_u411  (
    .a({\t/a/ID_rs1 [0],_al_u407_o}),
    .b({\t/a/ID_rs1 [1],_al_u408_o}),
    .c({\t/a/regfile/regfile$4$ [9],_al_u409_o}),
    .d({\t/a/regfile/regfile$5$ [9],_al_u410_o}),
    .e({open_n16182,\t/a/ID_rs1 [2]}),
    .f({_al_u344_o,_al_u411_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u353|t/a/regfile/reg0_b393  (
    .a({_al_u348_o,_al_u349_o}),
    .b({_al_u350_o,\t/a/ID_rs1 [0]}),
    .c({_al_u352_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [9]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [9]}),
    .mi({open_n16204,\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({_al_u353_o,_al_u350_o}),
    .q({open_n16219,\t/a/regfile/regfile$12$ [9]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u355|_al_u1085  (
    .a({\t/a/ID_rs1 [0],_al_u1081_o}),
    .b({\t/a/ID_rs1 [1],_al_u1082_o}),
    .c({\t/a/regfile/regfile$4$ [8],_al_u1083_o}),
    .d({\t/a/regfile/regfile$5$ [8],_al_u1084_o}),
    .e({open_n16222,\t/a/ID_rs2 [2]}),
    .f({_al_u355_o,_al_u1085_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u364|t/a/regfile/reg0_b392  (
    .a({_al_u359_o,_al_u360_o}),
    .b({_al_u361_o,\t/a/ID_rs1 [0]}),
    .c({_al_u363_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [8]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [8]}),
    .mi({open_n16244,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u364_o,_al_u361_o}),
    .q({open_n16259,\t/a/regfile/regfile$12$ [8]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u369|_al_u684  (
    .a({_al_u365_o,_al_u680_o}),
    .b({_al_u366_o,_al_u681_o}),
    .c({_al_u367_o,_al_u682_o}),
    .d({_al_u368_o,_al_u683_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .f({_al_u369_o,_al_u684_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u374|t/a/regfile/reg0_b904  (
    .a({_al_u369_o,_al_u370_o}),
    .b({_al_u371_o,\t/a/ID_rs1 [0]}),
    .c({_al_u373_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [8]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [8]}),
    .mi({open_n16283,\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u374_o,_al_u371_o}),
    .q({open_n16298,\t/a/regfile/regfile$28$ [8]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u380 (
    .a({_al_u376_o,_al_u376_o}),
    .b({_al_u377_o,_al_u377_o}),
    .c({_al_u378_o,_al_u378_o}),
    .d({_al_u379_o,_al_u379_o}),
    .mi({open_n16311,\t/a/ID_rs1 [2]}),
    .fx({open_n16316,_al_u380_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u385|t/a/regfile/reg0_b647  (
    .a({_al_u380_o,_al_u381_o}),
    .b({_al_u382_o,\t/a/ID_rs1 [0]}),
    .c({_al_u384_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [7]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [7]}),
    .mi({open_n16320,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({_al_u385_o,_al_u382_o}),
    .q({open_n16335,\t/a/regfile/regfile$20$ [7]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b0000010010001100),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000010010001100),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u386|_al_u1093  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$4$ [7],\t/a/regfile/regfile$6$ [7]}),
    .d({\t/a/regfile/regfile$5$ [7],\t/a/regfile/regfile$7$ [7]}),
    .f({_al_u386_o,_al_u1093_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u390 (
    .a({_al_u386_o,_al_u386_o}),
    .b({_al_u387_o,_al_u387_o}),
    .c({_al_u388_o,_al_u388_o}),
    .d({_al_u389_o,_al_u389_o}),
    .mi({open_n16372,\t/a/ID_rs1 [2]}),
    .fx({open_n16377,_al_u390_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u395|t/a/regfile/reg0_b391  (
    .a({_al_u390_o,_al_u391_o}),
    .b({_al_u392_o,\t/a/ID_rs1 [0]}),
    .c({_al_u394_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [7]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [7]}),
    .mi({open_n16381,\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({_al_u395_o,_al_u392_o}),
    .q({open_n16396,\t/a/regfile/regfile$12$ [7]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u397|_al_u401  (
    .a({\t/a/ID_rs1 [0],_al_u397_o}),
    .b({\t/a/ID_rs1 [1],_al_u398_o}),
    .c({\t/a/regfile/regfile$4$ [6],_al_u399_o}),
    .d({\t/a/regfile/regfile$5$ [6],_al_u400_o}),
    .e({open_n16399,\t/a/ID_rs1 [2]}),
    .f({_al_u397_o,_al_u401_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u406|t/a/regfile/reg0_b390  (
    .a({_al_u401_o,_al_u402_o}),
    .b({_al_u403_o,\t/a/ID_rs1 [0]}),
    .c({_al_u405_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [6]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [6]}),
    .mi({open_n16421,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u406_o,_al_u403_o}),
    .q({open_n16436,\t/a/regfile/regfile$12$ [6]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u416|t/a/regfile/reg0_b902  (
    .a({_al_u411_o,_al_u412_o}),
    .b({_al_u413_o,\t/a/ID_rs1 [0]}),
    .c({_al_u415_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [6]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [6]}),
    .mi({open_n16438,\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u416_o,_al_u413_o}),
    .q({open_n16453,\t/a/regfile/regfile$28$ [6]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u422 (
    .a({_al_u418_o,_al_u418_o}),
    .b({_al_u419_o,_al_u419_o}),
    .c({_al_u420_o,_al_u420_o}),
    .d({_al_u421_o,_al_u421_o}),
    .mi({open_n16466,\t/a/ID_rs1 [2]}),
    .fx({open_n16471,_al_u422_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u427|t/a/regfile/reg0_b389  (
    .a({_al_u422_o,_al_u423_o}),
    .b({_al_u424_o,\t/a/ID_rs1 [0]}),
    .c({_al_u426_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [5]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [5]}),
    .mi({open_n16475,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u427_o,_al_u424_o}),
    .q({open_n16490,\t/a/regfile/regfile$12$ [5]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u432|_al_u621  (
    .a({_al_u428_o,_al_u617_o}),
    .b({_al_u429_o,_al_u618_o}),
    .c({_al_u430_o,_al_u619_o}),
    .d({_al_u431_o,_al_u620_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .f({_al_u432_o,_al_u621_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u437|t/a/regfile/reg0_b901  (
    .a({_al_u432_o,_al_u433_o}),
    .b({_al_u434_o,\t/a/ID_rs1 [0]}),
    .c({_al_u436_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [5]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [5]}),
    .mi({open_n16514,\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u437_o,_al_u434_o}),
    .q({open_n16529,\t/a/regfile/regfile$28$ [5]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u443 (
    .a({_al_u439_o,_al_u439_o}),
    .b({_al_u440_o,_al_u440_o}),
    .c({_al_u441_o,_al_u441_o}),
    .d({_al_u442_o,_al_u442_o}),
    .mi({open_n16542,\t/a/ID_rs1 [2]}),
    .fx({open_n16547,_al_u443_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u448|t/a/regfile/reg0_b644  (
    .a({_al_u443_o,_al_u444_o}),
    .b({_al_u445_o,\t/a/ID_rs1 [0]}),
    .c({_al_u447_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [4]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [4]}),
    .mi({open_n16551,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u448_o,_al_u445_o}),
    .q({open_n16566,\t/a/regfile/regfile$20$ [4]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u449|_al_u453  (
    .a({\t/a/ID_rs1 [0],_al_u449_o}),
    .b({\t/a/ID_rs1 [1],_al_u450_o}),
    .c({\t/a/regfile/regfile$4$ [4],_al_u451_o}),
    .d({\t/a/regfile/regfile$5$ [4],_al_u452_o}),
    .e({open_n16569,\t/a/ID_rs1 [2]}),
    .f({_al_u449_o,_al_u453_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u450|_al_u1159  (
    .a({\t/a/ID_rs1 [0],_al_u1155_o}),
    .b({\t/a/ID_rs1 [1],_al_u1156_o}),
    .c({\t/a/regfile/regfile$6$ [4],_al_u1157_o}),
    .d({\t/a/regfile/regfile$7$ [4],_al_u1158_o}),
    .e({open_n16592,\t/a/ID_rs2 [2]}),
    .f({_al_u450_o,_al_u1159_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u458|t/a/regfile/reg0_b388  (
    .a({_al_u453_o,_al_u454_o}),
    .b({_al_u455_o,\t/a/ID_rs1 [0]}),
    .c({_al_u457_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [4]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [4]}),
    .mi({open_n16614,\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u458_o,_al_u455_o}),
    .q({open_n16629,\t/a/regfile/regfile$12$ [4]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u460|_al_u464  (
    .a({\t/a/ID_rs1 [0],_al_u460_o}),
    .b({\t/a/ID_rs1 [1],_al_u461_o}),
    .c({\t/a/regfile/regfile$4$ [3],_al_u462_o}),
    .d({\t/a/regfile/regfile$5$ [3],_al_u463_o}),
    .e({open_n16632,\t/a/ID_rs1 [2]}),
    .f({_al_u460_o,_al_u464_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u469|t/a/regfile/reg0_b387  (
    .a({_al_u464_o,_al_u465_o}),
    .b({_al_u466_o,\t/a/ID_rs1 [0]}),
    .c({_al_u468_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [3]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [3]}),
    .mi({open_n16654,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u469_o,_al_u466_o}),
    .q({open_n16669,\t/a/regfile/regfile$12$ [3]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u474|_al_u579  (
    .a({_al_u470_o,_al_u575_o}),
    .b({_al_u471_o,_al_u576_o}),
    .c({_al_u472_o,_al_u577_o}),
    .d({_al_u473_o,_al_u578_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .f({_al_u474_o,_al_u579_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u479|t/a/regfile/reg0_b899  (
    .a({_al_u474_o,_al_u475_o}),
    .b({_al_u476_o,\t/a/ID_rs1 [0]}),
    .c({_al_u478_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [3]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [3]}),
    .mi({open_n16693,\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u479_o,_al_u476_o}),
    .q({open_n16708,\t/a/regfile/regfile$28$ [3]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u485 (
    .a({_al_u481_o,_al_u481_o}),
    .b({_al_u482_o,_al_u482_o}),
    .c({_al_u483_o,_al_u483_o}),
    .d({_al_u484_o,_al_u484_o}),
    .mi({open_n16721,\t/a/ID_rs1 [2]}),
    .fx({open_n16726,_al_u485_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u490|t/a/regfile/reg0_b671  (
    .a({_al_u485_o,_al_u486_o}),
    .b({_al_u487_o,\t/a/ID_rs1 [0]}),
    .c({_al_u489_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [31]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [31]}),
    .mi({open_n16730,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u490_o,_al_u487_o}),
    .q({open_n16745,\t/a/regfile/regfile$20$ [31]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u495 (
    .a({_al_u491_o,_al_u491_o}),
    .b({_al_u492_o,_al_u492_o}),
    .c({_al_u493_o,_al_u493_o}),
    .d({_al_u494_o,_al_u494_o}),
    .mi({open_n16758,\t/a/ID_rs1 [2]}),
    .fx({open_n16763,_al_u495_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u500|t/a/regfile/reg0_b415  (
    .a({_al_u495_o,_al_u496_o}),
    .b({_al_u497_o,\t/a/ID_rs1 [0]}),
    .c({_al_u499_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [31]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [31]}),
    .mi({open_n16767,\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u500_o,_al_u497_o}),
    .q({open_n16782,\t/a/regfile/regfile$12$ [31]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u502|_al_u506  (
    .a({\t/a/ID_rs1 [0],_al_u502_o}),
    .b({\t/a/ID_rs1 [1],_al_u503_o}),
    .c({\t/a/regfile/regfile$4$ [30],_al_u504_o}),
    .d({\t/a/regfile/regfile$5$ [30],_al_u505_o}),
    .e({open_n16785,\t/a/ID_rs1 [2]}),
    .f({_al_u502_o,_al_u506_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u511|t/a/regfile/reg0_b414  (
    .a({_al_u506_o,_al_u507_o}),
    .b({_al_u508_o,\t/a/ID_rs1 [0]}),
    .c({_al_u510_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [30]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [30]}),
    .mi({open_n16807,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u511_o,_al_u508_o}),
    .q({open_n16822,\t/a/regfile/regfile$12$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u516|_al_u768  (
    .a({_al_u512_o,_al_u764_o}),
    .b({_al_u513_o,_al_u765_o}),
    .c({_al_u514_o,_al_u766_o}),
    .d({_al_u515_o,_al_u767_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .f({_al_u516_o,_al_u768_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u521|t/a/regfile/reg0_b926  (
    .a({_al_u516_o,_al_u517_o}),
    .b({_al_u518_o,\t/a/ID_rs1 [0]}),
    .c({_al_u520_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [30]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [30]}),
    .mi({open_n16846,\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u521_o,_al_u518_o}),
    .q({open_n16861,\t/a/regfile/regfile$28$ [30]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u523|_al_u527  (
    .a({\t/a/ID_rs1 [0],_al_u523_o}),
    .b({\t/a/ID_rs1 [1],_al_u524_o}),
    .c({\t/a/regfile/regfile$4$ [2],_al_u525_o}),
    .d({\t/a/regfile/regfile$5$ [2],_al_u526_o}),
    .e({open_n16864,\t/a/ID_rs1 [2]}),
    .f({_al_u523_o,_al_u527_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u532|t/a/regfile/reg0_b386  (
    .a({_al_u527_o,_al_u528_o}),
    .b({_al_u529_o,\t/a/ID_rs1 [0]}),
    .c({_al_u531_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [2]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [2]}),
    .mi({open_n16886,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u532_o,_al_u529_o}),
    .q({open_n16901,\t/a/regfile/regfile$12$ [2]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u537 (
    .a({_al_u533_o,_al_u533_o}),
    .b({_al_u534_o,_al_u534_o}),
    .c({_al_u535_o,_al_u535_o}),
    .d({_al_u536_o,_al_u536_o}),
    .mi({open_n16914,\t/a/ID_rs1 [2]}),
    .fx({open_n16919,_al_u537_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u542|t/a/regfile/reg0_b898  (
    .a({_al_u537_o,_al_u538_o}),
    .b({_al_u539_o,\t/a/ID_rs1 [0]}),
    .c({_al_u541_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [2]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [2]}),
    .mi({open_n16923,\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u542_o,_al_u539_o}),
    .q({open_n16938,\t/a/regfile/regfile$28$ [2]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u548 (
    .a({_al_u544_o,_al_u544_o}),
    .b({_al_u545_o,_al_u545_o}),
    .c({_al_u546_o,_al_u546_o}),
    .d({_al_u547_o,_al_u547_o}),
    .mi({open_n16951,\t/a/ID_rs1 [2]}),
    .fx({open_n16956,_al_u548_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u553|t/a/regfile/reg0_b669  (
    .a({_al_u548_o,_al_u549_o}),
    .b({_al_u550_o,\t/a/ID_rs1 [0]}),
    .c({_al_u552_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [29]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [29]}),
    .mi({open_n16960,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u553_o,_al_u550_o}),
    .q({open_n16975,\t/a/regfile/regfile$20$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u554|_al_u1260  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$4$ [29],\t/a/regfile/regfile$4$ [29]}),
    .d({\t/a/regfile/regfile$5$ [29],\t/a/regfile/regfile$5$ [29]}),
    .f({_al_u554_o,_al_u1260_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u558|_al_u810  (
    .a({_al_u554_o,_al_u806_o}),
    .b({_al_u555_o,_al_u807_o}),
    .c({_al_u556_o,_al_u808_o}),
    .d({_al_u557_o,_al_u809_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .f({_al_u558_o,_al_u810_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u563|t/a/regfile/reg0_b413  (
    .a({_al_u558_o,_al_u559_o}),
    .b({_al_u560_o,\t/a/ID_rs1 [0]}),
    .c({_al_u562_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [29]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [29]}),
    .mi({open_n17023,\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u563_o,_al_u560_o}),
    .q({open_n17038,\t/a/regfile/regfile$12$ [29]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u565|_al_u569  (
    .a({\t/a/ID_rs1 [0],_al_u565_o}),
    .b({\t/a/ID_rs1 [1],_al_u566_o}),
    .c({\t/a/regfile/regfile$4$ [28],_al_u567_o}),
    .d({\t/a/regfile/regfile$5$ [28],_al_u568_o}),
    .e({open_n17041,\t/a/ID_rs1 [2]}),
    .f({_al_u565_o,_al_u569_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u574|t/a/regfile/reg0_b412  (
    .a({_al_u569_o,_al_u570_o}),
    .b({_al_u571_o,\t/a/ID_rs1 [0]}),
    .c({_al_u573_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [28]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [28]}),
    .mi({open_n17063,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u574_o,_al_u571_o}),
    .q({open_n17078,\t/a/regfile/regfile$12$ [28]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u584|t/a/regfile/reg0_b924  (
    .a({_al_u579_o,_al_u580_o}),
    .b({_al_u581_o,\t/a/ID_rs1 [0]}),
    .c({_al_u583_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [28]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [28]}),
    .mi({open_n17080,\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u584_o,_al_u581_o}),
    .q({open_n17095,\t/a/regfile/regfile$28$ [28]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u590|_al_u800  (
    .a({_al_u586_o,_al_u796_o}),
    .b({_al_u587_o,_al_u797_o}),
    .c({_al_u588_o,_al_u798_o}),
    .d({_al_u589_o,_al_u799_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .f({_al_u590_o,_al_u800_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u595|t/a/regfile/reg0_b667  (
    .a({_al_u590_o,_al_u591_o}),
    .b({_al_u592_o,\t/a/ID_rs1 [0]}),
    .c({_al_u594_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [27]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [27]}),
    .mi({open_n17119,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u595_o,_al_u592_o}),
    .q({open_n17134,\t/a/regfile/regfile$20$ [27]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u600 (
    .a({_al_u596_o,_al_u596_o}),
    .b({_al_u597_o,_al_u597_o}),
    .c({_al_u598_o,_al_u598_o}),
    .d({_al_u599_o,_al_u599_o}),
    .mi({open_n17147,\t/a/ID_rs1 [2]}),
    .fx({open_n17152,_al_u600_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u605|t/a/regfile/reg0_b411  (
    .a({_al_u600_o,_al_u601_o}),
    .b({_al_u602_o,\t/a/ID_rs1 [0]}),
    .c({_al_u604_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [27]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [27]}),
    .mi({open_n17156,\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u605_o,_al_u602_o}),
    .q({open_n17171,\t/a/regfile/regfile$12$ [27]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u607|_al_u1333  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$4$ [26],\t/a/regfile/regfile$4$ [26]}),
    .d({\t/a/regfile/regfile$5$ [26],\t/a/regfile/regfile$5$ [26]}),
    .f({_al_u607_o,_al_u1333_o}));
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u611 (
    .a({_al_u607_o,_al_u607_o}),
    .b({_al_u608_o,_al_u608_o}),
    .c({_al_u609_o,_al_u609_o}),
    .d({_al_u610_o,_al_u610_o}),
    .mi({open_n17208,\t/a/ID_rs1 [2]}),
    .fx({open_n17213,_al_u611_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u616|t/a/regfile/reg0_b410  (
    .a({_al_u611_o,_al_u612_o}),
    .b({_al_u613_o,\t/a/ID_rs1 [0]}),
    .c({_al_u615_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [26]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [26]}),
    .mi({open_n17217,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u616_o,_al_u613_o}),
    .q({open_n17232,\t/a/regfile/regfile$12$ [26]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u626|t/a/regfile/reg0_b922  (
    .a({_al_u621_o,_al_u622_o}),
    .b({_al_u623_o,\t/a/ID_rs1 [0]}),
    .c({_al_u625_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [26]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [26]}),
    .mi({open_n17234,\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u626_o,_al_u623_o}),
    .q({open_n17249,\t/a/regfile/regfile$28$ [26]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u628|_al_u632  (
    .a({\t/a/ID_rs1 [0],_al_u628_o}),
    .b({\t/a/ID_rs1 [1],_al_u629_o}),
    .c({\t/a/regfile/regfile$4$ [25],_al_u630_o}),
    .d({\t/a/regfile/regfile$5$ [25],_al_u631_o}),
    .e({open_n17252,\t/a/ID_rs1 [2]}),
    .f({_al_u628_o,_al_u632_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u637|t/a/regfile/reg0_b409  (
    .a({_al_u632_o,_al_u633_o}),
    .b({_al_u634_o,\t/a/ID_rs1 [0]}),
    .c({_al_u636_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [25]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [25]}),
    .mi({open_n17274,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u637_o,_al_u634_o}),
    .q({open_n17289,\t/a/regfile/regfile$12$ [25]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u642 (
    .a({_al_u638_o,_al_u638_o}),
    .b({_al_u639_o,_al_u639_o}),
    .c({_al_u640_o,_al_u640_o}),
    .d({_al_u641_o,_al_u641_o}),
    .mi({open_n17302,\t/a/ID_rs1 [2]}),
    .fx({open_n17307,_al_u642_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u647|t/a/regfile/reg0_b921  (
    .a({_al_u642_o,_al_u643_o}),
    .b({_al_u644_o,\t/a/ID_rs1 [0]}),
    .c({_al_u646_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [25]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [25]}),
    .mi({open_n17311,\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u647_o,_al_u644_o}),
    .q({open_n17326,\t/a/regfile/regfile$28$ [25]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u653|_al_u957  (
    .a({_al_u649_o,_al_u953_o}),
    .b({_al_u650_o,_al_u954_o}),
    .c({_al_u651_o,_al_u955_o}),
    .d({_al_u652_o,_al_u956_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .f({_al_u653_o,_al_u957_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u658|t/a/regfile/reg0_b408  (
    .a({_al_u653_o,_al_u654_o}),
    .b({_al_u655_o,\t/a/ID_rs1 [0]}),
    .c({_al_u657_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [24]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [24]}),
    .mi({open_n17350,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u658_o,_al_u655_o}),
    .q({open_n17365,\t/a/regfile/regfile$12$ [24]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u663 (
    .a({_al_u659_o,_al_u659_o}),
    .b({_al_u660_o,_al_u660_o}),
    .c({_al_u661_o,_al_u661_o}),
    .d({_al_u662_o,_al_u662_o}),
    .mi({open_n17378,\t/a/ID_rs1 [2]}),
    .fx({open_n17383,_al_u663_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u668|t/a/regfile/reg0_b920  (
    .a({_al_u663_o,_al_u664_o}),
    .b({_al_u665_o,\t/a/ID_rs1 [0]}),
    .c({_al_u667_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [24]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [24]}),
    .mi({open_n17387,\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u668_o,_al_u665_o}),
    .q({open_n17402,\t/a/regfile/regfile$28$ [24]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u670|_al_u674  (
    .a({\t/a/ID_rs1 [0],_al_u670_o}),
    .b({\t/a/ID_rs1 [1],_al_u671_o}),
    .c({\t/a/regfile/regfile$4$ [23],_al_u672_o}),
    .d({\t/a/regfile/regfile$5$ [23],_al_u673_o}),
    .e({open_n17405,\t/a/ID_rs1 [2]}),
    .f({_al_u670_o,_al_u674_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u679|t/a/regfile/reg0_b407  (
    .a({_al_u674_o,_al_u675_o}),
    .b({_al_u676_o,\t/a/ID_rs1 [0]}),
    .c({_al_u678_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [23]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [23]}),
    .mi({open_n17427,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u679_o,_al_u676_o}),
    .q({open_n17442,\t/a/regfile/regfile$12$ [23]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u689|t/a/regfile/reg0_b919  (
    .a({_al_u684_o,_al_u685_o}),
    .b({_al_u686_o,\t/a/ID_rs1 [0]}),
    .c({_al_u688_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [23]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [23]}),
    .mi({open_n17444,\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u689_o,_al_u686_o}),
    .q({open_n17459,\t/a/regfile/regfile$28$ [23]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u695|_al_u947  (
    .a({_al_u691_o,_al_u943_o}),
    .b({_al_u692_o,_al_u944_o}),
    .c({_al_u693_o,_al_u945_o}),
    .d({_al_u694_o,_al_u946_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .f({_al_u695_o,_al_u947_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u700|t/a/regfile/reg0_b662  (
    .a({_al_u695_o,_al_u696_o}),
    .b({_al_u697_o,\t/a/ID_rs1 [0]}),
    .c({_al_u699_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [22]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [22]}),
    .mi({open_n17483,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u700_o,_al_u697_o}),
    .q({open_n17498,\t/a/regfile/regfile$20$ [22]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u701|t/a/regfile/reg0_b182  (
    .a({\t/a/ID_rs1 [0],_al_u1853_o}),
    .b({\t/a/ID_rs1 [1],\t/a/alu_A_select [1]}),
    .c({\t/a/regfile/regfile$4$ [22],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [22],\t/a/reg_writedat [22]}),
    .mi({open_n17509,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u701_o,\t/a/aluin/sel0_b22/B0 }),
    .q({open_n17513,\t/a/regfile/regfile$5$ [22]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u705|_al_u1411  (
    .a({_al_u701_o,_al_u1407_o}),
    .b({_al_u702_o,_al_u1408_o}),
    .c({_al_u703_o,_al_u1409_o}),
    .d({_al_u704_o,_al_u1410_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs2 [2]}),
    .f({_al_u705_o,_al_u1411_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u710|t/a/regfile/reg0_b406  (
    .a({_al_u705_o,_al_u706_o}),
    .b({_al_u707_o,\t/a/ID_rs1 [0]}),
    .c({_al_u709_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [22]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [22]}),
    .mi({open_n17537,\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u710_o,_al_u707_o}),
    .q({open_n17552,\t/a/regfile/regfile$12$ [22]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u712|t/a/regfile/reg0_b181  (
    .a({\t/a/ID_rs1 [0],_al_u1856_o}),
    .b({\t/a/ID_rs1 [1],\t/a/alu_A_select [1]}),
    .c({\t/a/regfile/regfile$4$ [21],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [21],\t/a/reg_writedat [21]}),
    .mi({open_n17563,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u712_o,\t/a/aluin/sel0_b21/B0 }),
    .q({open_n17567,\t/a/regfile/regfile$5$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u716 (
    .a({_al_u712_o,_al_u712_o}),
    .b({_al_u713_o,_al_u713_o}),
    .c({_al_u714_o,_al_u714_o}),
    .d({_al_u715_o,_al_u715_o}),
    .mi({open_n17580,\t/a/ID_rs1 [2]}),
    .fx({open_n17585,_al_u716_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u721|t/a/regfile/reg0_b405  (
    .a({_al_u716_o,_al_u717_o}),
    .b({_al_u718_o,\t/a/ID_rs1 [0]}),
    .c({_al_u720_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [21]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [21]}),
    .mi({open_n17589,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u721_o,_al_u718_o}),
    .q({open_n17604,\t/a/regfile/regfile$12$ [21]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u726 (
    .a({_al_u722_o,_al_u722_o}),
    .b({_al_u723_o,_al_u723_o}),
    .c({_al_u724_o,_al_u724_o}),
    .d({_al_u725_o,_al_u725_o}),
    .mi({open_n17617,\t/a/ID_rs1 [2]}),
    .fx({open_n17622,_al_u726_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u731|t/a/regfile/reg0_b917  (
    .a({_al_u726_o,_al_u727_o}),
    .b({_al_u728_o,\t/a/ID_rs1 [0]}),
    .c({_al_u730_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [21]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [21]}),
    .mi({open_n17626,\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u731_o,_al_u728_o}),
    .q({open_n17641,\t/a/regfile/regfile$28$ [21]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u737|_al_u905  (
    .a({_al_u733_o,_al_u901_o}),
    .b({_al_u734_o,_al_u902_o}),
    .c({_al_u735_o,_al_u903_o}),
    .d({_al_u736_o,_al_u904_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .f({_al_u737_o,_al_u905_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u742|t/a/regfile/reg0_b660  (
    .a({_al_u737_o,_al_u738_o}),
    .b({_al_u739_o,\t/a/ID_rs1 [0]}),
    .c({_al_u741_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [20]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [20]}),
    .mi({open_n17665,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u742_o,_al_u739_o}),
    .q({open_n17680,\t/a/regfile/regfile$20$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u747|_al_u863  (
    .a({_al_u743_o,_al_u859_o}),
    .b({_al_u744_o,_al_u860_o}),
    .c({_al_u745_o,_al_u861_o}),
    .d({_al_u746_o,_al_u862_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .f({_al_u747_o,_al_u863_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u752|t/a/regfile/reg0_b404  (
    .a({_al_u747_o,_al_u748_o}),
    .b({_al_u749_o,\t/a/ID_rs1 [0]}),
    .c({_al_u751_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [20]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [20]}),
    .mi({open_n17704,\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u752_o,_al_u749_o}),
    .q({open_n17719,\t/a/regfile/regfile$12$ [20]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u754|_al_u758  (
    .a({\t/a/ID_rs1 [0],_al_u754_o}),
    .b({\t/a/ID_rs1 [1],_al_u755_o}),
    .c({\t/a/regfile/regfile$4$ [1],_al_u756_o}),
    .d({\t/a/regfile/regfile$5$ [1],_al_u757_o}),
    .e({open_n17722,\t/a/ID_rs1 [2]}),
    .f({_al_u754_o,_al_u758_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u763|t/a/regfile/reg0_b385  (
    .a({_al_u758_o,_al_u759_o}),
    .b({_al_u760_o,\t/a/ID_rs1 [0]}),
    .c({_al_u762_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [1]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [1]}),
    .mi({open_n17744,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u763_o,_al_u760_o}),
    .q({open_n17759,\t/a/regfile/regfile$12$ [1]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u773|t/a/regfile/reg0_b897  (
    .a({_al_u768_o,_al_u769_o}),
    .b({_al_u770_o,\t/a/ID_rs1 [0]}),
    .c({_al_u772_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [1]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [1]}),
    .mi({open_n17761,\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u773_o,_al_u770_o}),
    .q({open_n17776,\t/a/regfile/regfile$28$ [1]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~A*~(~D*B))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*~A*~(~D*B))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101000000010000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u775|t/a/regfile/reg0_b179  (
    .a({\t/a/ID_rs1 [0],_al_u1865_o}),
    .b({\t/a/ID_rs1 [1],\t/a/alu_A_select [1]}),
    .c({\t/a/regfile/regfile$4$ [19],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [19],\t/a/reg_writedat [19]}),
    .mi({open_n17780,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u775_o,\t/a/aluin/sel0_b19/B0 }),
    .q({open_n17795,\t/a/regfile/regfile$5$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u779 (
    .a({_al_u775_o,_al_u775_o}),
    .b({_al_u776_o,_al_u776_o}),
    .c({_al_u777_o,_al_u777_o}),
    .d({_al_u778_o,_al_u778_o}),
    .mi({open_n17808,\t/a/ID_rs1 [2]}),
    .fx({open_n17813,_al_u779_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u784|t/a/regfile/reg0_b403  (
    .a({_al_u779_o,_al_u780_o}),
    .b({_al_u781_o,\t/a/ID_rs1 [0]}),
    .c({_al_u783_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [19]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [19]}),
    .mi({open_n17817,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u784_o,_al_u781_o}),
    .q({open_n17832,\t/a/regfile/regfile$12$ [19]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u789 (
    .a({_al_u785_o,_al_u785_o}),
    .b({_al_u786_o,_al_u786_o}),
    .c({_al_u787_o,_al_u787_o}),
    .d({_al_u788_o,_al_u788_o}),
    .mi({open_n17845,\t/a/ID_rs1 [2]}),
    .fx({open_n17850,_al_u789_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u794|t/a/regfile/reg0_b915  (
    .a({_al_u789_o,_al_u790_o}),
    .b({_al_u791_o,\t/a/ID_rs1 [0]}),
    .c({_al_u793_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [19]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [19]}),
    .mi({open_n17854,\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u794_o,_al_u791_o}),
    .q({open_n17869,\t/a/regfile/regfile$28$ [19]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u805|t/a/regfile/reg0_b658  (
    .a({_al_u800_o,_al_u801_o}),
    .b({_al_u802_o,\t/a/ID_rs1 [0]}),
    .c({_al_u804_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [18]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [18]}),
    .mi({open_n17871,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u805_o,_al_u802_o}),
    .q({open_n17886,\t/a/regfile/regfile$20$ [18]}));  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u806|t/a/regfile/reg0_b178  (
    .a({\t/a/ID_rs1 [0],_al_u1868_o}),
    .b({\t/a/ID_rs1 [1],\t/a/alu_A_select [1]}),
    .c({\t/a/regfile/regfile$4$ [18],\t/a/aluin/n5_lutinv }),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [18],\t/a/reg_writedat [18]}),
    .mi({open_n17897,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u806_o,\t/a/aluin/sel0_b18/B0 }),
    .q({open_n17901,\t/a/regfile/regfile$5$ [18]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u815|t/a/regfile/reg0_b402  (
    .a({_al_u810_o,_al_u811_o}),
    .b({_al_u812_o,\t/a/ID_rs1 [0]}),
    .c({_al_u814_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [18]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [18]}),
    .mi({open_n17903,\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u815_o,_al_u812_o}),
    .q({open_n17918,\t/a/regfile/regfile$12$ [18]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u821 (
    .a({_al_u817_o,_al_u817_o}),
    .b({_al_u818_o,_al_u818_o}),
    .c({_al_u819_o,_al_u819_o}),
    .d({_al_u820_o,_al_u820_o}),
    .mi({open_n17931,\t/a/ID_rs1 [2]}),
    .fx({open_n17936,_al_u821_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u826|t/a/regfile/reg0_b401  (
    .a({_al_u821_o,_al_u822_o}),
    .b({_al_u823_o,\t/a/ID_rs1 [0]}),
    .c({_al_u825_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [17]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [17]}),
    .mi({open_n17940,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u826_o,_al_u823_o}),
    .q({open_n17955,\t/a/regfile/regfile$12$ [17]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u831|_al_u873  (
    .a({_al_u827_o,_al_u869_o}),
    .b({_al_u828_o,_al_u870_o}),
    .c({_al_u829_o,_al_u871_o}),
    .d({_al_u830_o,_al_u872_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .f({_al_u831_o,_al_u873_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u836|t/a/regfile/reg0_b913  (
    .a({_al_u831_o,_al_u832_o}),
    .b({_al_u833_o,\t/a/ID_rs1 [0]}),
    .c({_al_u835_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [17]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [17]}),
    .mi({open_n17979,\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u836_o,_al_u833_o}),
    .q({open_n17994,\t/a/regfile/regfile$28$ [17]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u842 (
    .a({_al_u838_o,_al_u838_o}),
    .b({_al_u839_o,_al_u839_o}),
    .c({_al_u840_o,_al_u840_o}),
    .d({_al_u841_o,_al_u841_o}),
    .mi({open_n18007,\t/a/ID_rs1 [2]}),
    .fx({open_n18012,_al_u842_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u847|t/a/regfile/reg0_b656  (
    .a({_al_u842_o,_al_u843_o}),
    .b({_al_u844_o,\t/a/ID_rs1 [0]}),
    .c({_al_u846_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [16]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [16]}),
    .mi({open_n18016,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u847_o,_al_u844_o}),
    .q({open_n18031,\t/a/regfile/regfile$20$ [16]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b1111111111110000),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b1110111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u852|_al_u1558  (
    .a({_al_u848_o,_al_u1554_o}),
    .b({_al_u849_o,_al_u1555_o}),
    .c({_al_u850_o,_al_u1556_o}),
    .d({_al_u851_o,_al_u1557_o}),
    .e({\t/a/ID_rs1 [2],\t/a/ID_rs2 [2]}),
    .f({_al_u852_o,_al_u1558_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u857|t/a/regfile/reg0_b400  (
    .a({_al_u852_o,_al_u853_o}),
    .b({_al_u854_o,\t/a/ID_rs1 [0]}),
    .c({_al_u856_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [16]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [16]}),
    .mi({open_n18055,\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u857_o,_al_u854_o}),
    .q({open_n18070,\t/a/regfile/regfile$12$ [16]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u868|t/a/regfile/reg0_b399  (
    .a({_al_u863_o,_al_u864_o}),
    .b({_al_u865_o,\t/a/ID_rs1 [0]}),
    .c({_al_u867_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [15]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [15]}),
    .mi({open_n18072,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u868_o,_al_u865_o}),
    .q({open_n18087,\t/a/regfile/regfile$12$ [15]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u878|t/a/regfile/reg0_b911  (
    .a({_al_u873_o,_al_u874_o}),
    .b({_al_u875_o,\t/a/ID_rs1 [0]}),
    .c({_al_u877_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [15]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [15]}),
    .mi({open_n18089,\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u878_o,_al_u875_o}),
    .q({open_n18104,\t/a/regfile/regfile$28$ [15]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u884 (
    .a({_al_u880_o,_al_u880_o}),
    .b({_al_u881_o,_al_u881_o}),
    .c({_al_u882_o,_al_u882_o}),
    .d({_al_u883_o,_al_u883_o}),
    .mi({open_n18117,\t/a/ID_rs1 [2]}),
    .fx({open_n18122,_al_u884_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u889|t/a/regfile/reg0_b398  (
    .a({_al_u884_o,_al_u885_o}),
    .b({_al_u886_o,\t/a/ID_rs1 [0]}),
    .c({_al_u888_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [14]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [14]}),
    .mi({open_n18126,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u889_o,_al_u886_o}),
    .q({open_n18141,\t/a/regfile/regfile$12$ [14]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u894 (
    .a({_al_u890_o,_al_u890_o}),
    .b({_al_u891_o,_al_u891_o}),
    .c({_al_u892_o,_al_u892_o}),
    .d({_al_u893_o,_al_u893_o}),
    .mi({open_n18154,\t/a/ID_rs1 [2]}),
    .fx({open_n18159,_al_u894_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u899|t/a/regfile/reg0_b910  (
    .a({_al_u894_o,_al_u895_o}),
    .b({_al_u896_o,\t/a/ID_rs1 [0]}),
    .c({_al_u898_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [14]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [14]}),
    .mi({open_n18163,\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u899_o,_al_u896_o}),
    .q({open_n18178,\t/a/regfile/regfile$28$ [14]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u910|t/a/regfile/reg0_b653  (
    .a({_al_u905_o,_al_u906_o}),
    .b({_al_u907_o,\t/a/ID_rs1 [0]}),
    .c({_al_u909_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [13]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [13]}),
    .mi({open_n18180,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u910_o,_al_u907_o}),
    .q({open_n18195,\t/a/regfile/regfile$20$ [13]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u920|t/a/regfile/reg0_b397  (
    .a({_al_u915_o,_al_u916_o}),
    .b({_al_u917_o,\t/a/ID_rs1 [0]}),
    .c({_al_u919_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [13]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [13]}),
    .mi({open_n18197,\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u920_o,_al_u917_o}),
    .q({open_n18212,\t/a/regfile/regfile$12$ [13]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u926 (
    .a({_al_u922_o,_al_u922_o}),
    .b({_al_u923_o,_al_u923_o}),
    .c({_al_u924_o,_al_u924_o}),
    .d({_al_u925_o,_al_u925_o}),
    .mi({open_n18225,\t/a/ID_rs1 [2]}),
    .fx({open_n18230,_al_u926_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u931|t/a/regfile/reg0_b396  (
    .a({_al_u926_o,_al_u927_o}),
    .b({_al_u928_o,\t/a/ID_rs1 [0]}),
    .c({_al_u930_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [12]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [12]}),
    .mi({open_n18234,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u931_o,_al_u928_o}),
    .q({open_n18249,\t/a/regfile/regfile$12$ [12]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u936 (
    .a({_al_u932_o,_al_u932_o}),
    .b({_al_u933_o,_al_u933_o}),
    .c({_al_u934_o,_al_u934_o}),
    .d({_al_u935_o,_al_u935_o}),
    .mi({open_n18262,\t/a/ID_rs1 [2]}),
    .fx({open_n18267,_al_u936_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u941|t/a/regfile/reg0_b908  (
    .a({_al_u936_o,_al_u937_o}),
    .b({_al_u938_o,\t/a/ID_rs1 [0]}),
    .c({_al_u940_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [12]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [12]}),
    .mi({open_n18271,\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u941_o,_al_u938_o}),
    .q({open_n18286,\t/a/regfile/regfile$28$ [12]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*((~C*~B)*~(A)*~(D)+(~C*~B)*A*~(D)+~((~C*~B))*A*D+(~C*~B)*A*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u952|t/a/regfile/reg0_b651  (
    .a({_al_u947_o,_al_u948_o}),
    .b({_al_u949_o,\t/a/ID_rs1 [0]}),
    .c({_al_u951_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$20$ [11]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$21$ [11]}),
    .mi({open_n18288,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u952_o,_al_u949_o}),
    .q({open_n18303,\t/a/regfile/regfile$20$ [11]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u962|t/a/regfile/reg0_b395  (
    .a({_al_u957_o,_al_u958_o}),
    .b({_al_u959_o,\t/a/ID_rs1 [0]}),
    .c({_al_u961_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [11]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [11]}),
    .mi({open_n18305,\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u962_o,_al_u959_o}),
    .q({open_n18320,\t/a/regfile/regfile$12$ [11]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u968 (
    .a({_al_u964_o,_al_u964_o}),
    .b({_al_u965_o,_al_u965_o}),
    .c({_al_u966_o,_al_u966_o}),
    .d({_al_u967_o,_al_u967_o}),
    .mi({open_n18333,\t/a/ID_rs1 [2]}),
    .fx({open_n18338,_al_u968_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u973|t/a/regfile/reg0_b394  (
    .a({_al_u968_o,_al_u969_o}),
    .b({_al_u970_o,\t/a/ID_rs1 [0]}),
    .c({_al_u972_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$12$ [10]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$13$ [10]}),
    .mi({open_n18342,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u973_o,_al_u970_o}),
    .q({open_n18357,\t/a/regfile/regfile$12$ [10]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUT1("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1110111011101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u978 (
    .a({_al_u974_o,_al_u974_o}),
    .b({_al_u975_o,_al_u975_o}),
    .c({_al_u976_o,_al_u976_o}),
    .d({_al_u977_o,_al_u977_o}),
    .mi({open_n18370,\t/a/ID_rs1 [2]}),
    .fx({open_n18375,_al_u978_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000001110101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u983|t/a/regfile/reg0_b906  (
    .a({_al_u978_o,_al_u979_o}),
    .b({_al_u980_o,\t/a/ID_rs1 [0]}),
    .c({_al_u982_o,\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$28$ [10]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$29$ [10]}),
    .mi({open_n18379,\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u983_o,_al_u980_o}),
    .q({open_n18394,\t/a/regfile/regfile$28$ [10]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*~C*~B*A)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~1*D*~C*~B*A)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u985|t/a/regfile/reg0_b128  (
    .a({\t/a/ID_rs1 [0],_al_u254_o}),
    .b({\t/a/ID_rs1 [1],\t/a/WB_rd [0]}),
    .c({\t/a/regfile/regfile$4$ [0],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$5$ [0],\t/a/WB_rd [2]}),
    .e({open_n18395,\t/a/WB_rd [3]}),
    .mi({open_n18397,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u985_o,\t/a/regfile/mux39_b128_sel_is_3_o }),
    .q({open_n18412,\t/a/regfile/regfile$4$ [0]}));  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*C*~B*A)"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~1*D*C*~B*A)"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u986|t/a/regfile/reg0_b192  (
    .a({\t/a/ID_rs1 [0],_al_u254_o}),
    .b({\t/a/ID_rs1 [1],\t/a/WB_rd [0]}),
    .c({\t/a/regfile/regfile$6$ [0],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [0],\t/a/WB_rd [2]}),
    .e({open_n18413,\t/a/WB_rd [3]}),
    .mi({open_n18415,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u986_o,\t/a/regfile/mux39_b192_sel_is_3_o }),
    .q({open_n18430,\t/a/regfile/regfile$6$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u987|_al_u989  (
    .a({\t/a/ID_rs1 [0],_al_u985_o}),
    .b({\t/a/ID_rs1 [1],_al_u986_o}),
    .c({\t/a/regfile/regfile$0$ [0],_al_u987_o}),
    .d({\t/a/regfile/regfile$1$ [0],_al_u988_o}),
    .e({open_n18433,\t/a/ID_rs1 [2]}),
    .f({_al_u987_o,_al_u989_o}));
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u988|t/a/regfile/reg0_b96  (
    .a({\t/a/ID_rs1 [0],_al_u2614_o}),
    .b({\t/a/ID_rs1 [1],_al_u2616_o}),
    .c({\t/a/regfile/regfile$2$ [0],\t/a/MEM_aludat [0]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$3$ [0],\t/a/reg_writedat [0]}),
    .mi({open_n18464,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u988_o,_al_u2760_o}),
    .q({open_n18468,\t/a/regfile/regfile$3$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u990|_al_u1706  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs2 [2]}),
    .d({\t/a/regfile/regfile$14$ [0],\t/a/regfile/regfile$14$ [0]}),
    .e({\t/a/regfile/regfile$15$ [0],\t/a/regfile/regfile$15$ [0]}),
    .f({_al_u990_o,_al_u1706_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*~B*A)"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(1*D*~C*~B*A)"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u991|t/a/regfile/reg0_b384  (
    .a({_al_u990_o,_al_u254_o}),
    .b({\t/a/ID_rs1 [0],\t/a/WB_rd [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$12$ [0],\t/a/WB_rd [2]}),
    .e({\t/a/regfile/regfile$13$ [0],\t/a/WB_rd [3]}),
    .mi({open_n18492,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u991_o,\t/a/regfile/mux39_b384_sel_is_3_o }),
    .q({open_n18507,\t/a/regfile/regfile$12$ [0]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUT1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .INIT_LUT0(16'b0000011100000011),
    .INIT_LUT1(16'b0000111100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u992 (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .d({\t/a/regfile/regfile$10$ [0],\t/a/regfile/regfile$10$ [0]}),
    .mi({open_n18520,\t/a/regfile/regfile$11$ [0]}),
    .fx({open_n18525,_al_u992_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*(A*~((~C*~B))*~(D)+A*(~C*~B)*~(D)+~(A)*(~C*~B)*D+A*(~C*~B)*D))"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000001110101010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u994|_al_u993  (
    .a({_al_u989_o,_al_u992_o}),
    .b({_al_u991_o,\t/a/ID_rs1 [0]}),
    .c({_al_u993_o,\t/a/ID_rs1 [1]}),
    .d({\t/a/ID_rs1 [3],\t/a/regfile/regfile$8$ [0]}),
    .e({\t/a/ID_rs1 [4],\t/a/regfile/regfile$9$ [0]}),
    .f({_al_u994_o,_al_u993_o}));
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*~C*~B*A)"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~1*D*~C*~B*A)"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u995|t/a/regfile/reg0_b640  (
    .a({\t/a/ID_rs1 [0],_al_u256_o}),
    .b({\t/a/ID_rs1 [1],\t/a/WB_rd [0]}),
    .c({\t/a/regfile/regfile$20$ [0],\t/a/WB_rd [1]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [0],\t/a/WB_rd [2]}),
    .e({open_n18550,\t/a/WB_rd [3]}),
    .mi({open_n18552,\t/a/reg_writedat [0]}),
    .sr(rst_pad),
    .f({_al_u995_o,\t/a/regfile/mux39_b640_sel_is_3_o }),
    .q({open_n18567,\t/a/regfile/regfile$20$ [0]}));  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("~((~D*~C)*~((~B*~A))*~(0)+(~D*~C)*(~B*~A)*~(0)+~((~D*~C))*(~B*~A)*0+(~D*~C)*(~B*~A)*0)"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("~((~D*~C)*~((~B*~A))*~(1)+(~D*~C)*(~B*~A)*~(1)+~((~D*~C))*(~B*~A)*1+(~D*~C)*(~B*~A)*1)"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b1110111011101110),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u996|_al_u999  (
    .a({\t/a/ID_rs1 [0],_al_u995_o}),
    .b({\t/a/ID_rs1 [1],_al_u996_o}),
    .c({\t/a/regfile/regfile$22$ [0],_al_u997_o}),
    .d({\t/a/regfile/regfile$23$ [0],_al_u998_o}),
    .e({open_n18570,\t/a/ID_rs1 [2]}),
    .f({_al_u996_o,_al_u999_o}));
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUTF0(16'b0000000100100011),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b0000000100100011),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u997|_al_u1713  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$16$ [0],\t/a/regfile/regfile$16$ [0]}),
    .d({\t/a/regfile/regfile$17$ [0],\t/a/regfile/regfile$17$ [0]}),
    .f({_al_u997_o,_al_u1713_o}));
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"))
    \_al_u998|_al_u1714  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$18$ [0],\t/a/regfile/regfile$18$ [0]}),
    .d({\t/a/regfile/regfile$19$ [0],\t/a/regfile/regfile$19$ [0]}),
    .f({_al_u998_o,_al_u1714_o}));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P138"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("RESET"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTRSTMUX("INV"),
    .OUTSCLKMUX("CLK"),
    .SRMODE("ASYNC"),
    .TSMUX("0"))
    led_n_reg_DO (
    .ce(n7),
    .do({open_n18682,open_n18683,open_n18684,o_data[0]}),
    .osclk(clock_pad),
    .rst(rst_pad),
    .opad(led));  // __top.v(63)
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_0|lt0_cin  (
    .a({addr[0],1'b0}),
    .b({1'b0,open_n18696}),
    .fco(lt0_c1));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_10|lt0_9  (
    .a(addr[10:9]),
    .b(2'b00),
    .fci(lt0_c9),
    .fco(lt0_c11));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_12|lt0_11  (
    .a(addr[12:11]),
    .b(2'b00),
    .fci(lt0_c11),
    .fco(lt0_c13));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_14|lt0_13  (
    .a(addr[14:13]),
    .b(2'b00),
    .fci(lt0_c13),
    .fco(lt0_c15));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_16|lt0_15  (
    .a(addr[16:15]),
    .b(2'b00),
    .fci(lt0_c15),
    .fco(lt0_c17));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_18|lt0_17  (
    .a(addr[18:17]),
    .b(2'b00),
    .fci(lt0_c17),
    .fco(lt0_c19));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_20|lt0_19  (
    .a(addr[20:19]),
    .b(2'b00),
    .fci(lt0_c19),
    .fco(lt0_c21));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_22|lt0_21  (
    .a(addr[22:21]),
    .b(2'b00),
    .fci(lt0_c21),
    .fco(lt0_c23));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_24|lt0_23  (
    .a(addr[24:23]),
    .b(2'b00),
    .fci(lt0_c23),
    .fco(lt0_c25));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_26|lt0_25  (
    .a(addr[26:25]),
    .b(2'b00),
    .fci(lt0_c25),
    .fco(lt0_c27));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_28|lt0_27  (
    .a(addr[28:27]),
    .b(2'b00),
    .fci(lt0_c27),
    .fco(lt0_c29));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_2|lt0_1  (
    .a(addr[2:1]),
    .b(2'b00),
    .fci(lt0_c1),
    .fco(lt0_c3));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_30|lt0_29  (
    .a(addr[30:29]),
    .b(2'b00),
    .fci(lt0_c29),
    .fco(lt0_c31));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_4|lt0_3  (
    .a(addr[4:3]),
    .b(2'b00),
    .fci(lt0_c3),
    .fco(lt0_c5));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_6|lt0_5  (
    .a(addr[6:5]),
    .b(2'b11),
    .fci(lt0_c5),
    .fco(lt0_c7));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_8|lt0_7  (
    .a(addr[8:7]),
    .b(2'b00),
    .fci(lt0_c7),
    .fco(lt0_c9));
  EG_PHY_MSLICE #(
    //.MACRO("lt0_0|lt0_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \lt0_cout|lt0_31  (
    .a({1'b0,addr[31]}),
    .b(2'b10),
    .fci(lt0_c31),
    .f({n0,open_n19100}));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c0_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c0_l  (
    .a({o_data[0],n2[0]}),
    .b({o_data[1],n2[1]}),
    .c({o_data[2],n2[2]}),
    .clk(clock_pad),
    .d({o_data[3],n2[3]}),
    .e({open_n19107,memwrite_cs}),
    .dpram_di(\m/dram_c0_di ),
    .dpram_mode(\m/dram_c0_mode ),
    .dpram_waddr(\m/dram_c0_waddr ),
    .dpram_wclk(\m/dram_c0_wclk ),
    .dpram_we(\m/dram_c0_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c0_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000110),
    .INIT_LUT1(16'b0000000000000110),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c0_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c0_di [1:0]),
    .dpram_mode(\m/dram_c0_mode ),
    .dpram_waddr(\m/dram_c0_waddr ),
    .dpram_wclk(\m/dram_c0_wclk ),
    .dpram_we(\m/dram_c0_we ),
    .sr(rst_pad),
    .f(i_data[1:0]),
    .q(\t/busarbitration/instruction [1:0]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c0_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c0_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c0_di [3:2]),
    .dpram_mode(\m/dram_c0_mode ),
    .dpram_waddr(\m/dram_c0_waddr ),
    .dpram_wclk(\m/dram_c0_wclk ),
    .dpram_we(\m/dram_c0_we ),
    .sr(rst_pad),
    .f(i_data[3:2]),
    .q(\t/busarbitration/instruction [3:2]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c1_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c1_l  (
    .a({o_data[4],n2[0]}),
    .b({o_data[5],n2[1]}),
    .c({o_data[6],n2[2]}),
    .clk(clock_pad),
    .d({o_data[7],n2[3]}),
    .e({open_n19132,memwrite_cs}),
    .dpram_di(\m/dram_c1_di ),
    .dpram_mode(\m/dram_c1_mode ),
    .dpram_waddr(\m/dram_c1_waddr ),
    .dpram_wclk(\m/dram_c1_wclk ),
    .dpram_we(\m/dram_c1_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c1_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000110),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c1_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c1_di [1:0]),
    .dpram_mode(\m/dram_c1_mode ),
    .dpram_waddr(\m/dram_c1_waddr ),
    .dpram_wclk(\m/dram_c1_wclk ),
    .dpram_we(\m/dram_c1_we ),
    .sr(rst_pad),
    .f(i_data[5:4]),
    .q(\t/busarbitration/instruction [5:4]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c1_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c1_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c1_di [3:2]),
    .dpram_mode(\m/dram_c1_mode ),
    .dpram_waddr(\m/dram_c1_waddr ),
    .dpram_wclk(\m/dram_c1_wclk ),
    .dpram_we(\m/dram_c1_we ),
    .sr(rst_pad),
    .f(i_data[7:6]),
    .q(\t/busarbitration/instruction [7:6]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c2_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c2_l  (
    .a({o_data[8],n2[0]}),
    .b({o_data[9],n2[1]}),
    .c({o_data[10],n2[2]}),
    .clk(clock_pad),
    .d({o_data[11],n2[3]}),
    .e({open_n19157,memwrite_cs}),
    .dpram_di(\m/dram_c2_di ),
    .dpram_mode(\m/dram_c2_mode ),
    .dpram_waddr(\m/dram_c2_waddr ),
    .dpram_wclk(\m/dram_c2_wclk ),
    .dpram_we(\m/dram_c2_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c2_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c2_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c2_di [1:0]),
    .dpram_mode(\m/dram_c2_mode ),
    .dpram_waddr(\m/dram_c2_waddr ),
    .dpram_wclk(\m/dram_c2_wclk ),
    .dpram_we(\m/dram_c2_we ),
    .sr(rst_pad),
    .f(i_data[9:8]),
    .q(\t/busarbitration/instruction [9:8]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c2_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c2_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c2_di [3:2]),
    .dpram_mode(\m/dram_c2_mode ),
    .dpram_waddr(\m/dram_c2_waddr ),
    .dpram_wclk(\m/dram_c2_wclk ),
    .dpram_we(\m/dram_c2_we ),
    .sr(rst_pad),
    .f(i_data[11:10]),
    .q(\t/busarbitration/instruction [11:10]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c3_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c3_l  (
    .a({o_data[12],n2[0]}),
    .b({o_data[13],n2[1]}),
    .c({o_data[14],n2[2]}),
    .clk(clock_pad),
    .d({o_data[15],n2[3]}),
    .e({open_n19182,memwrite_cs}),
    .dpram_di(\m/dram_c3_di ),
    .dpram_mode(\m/dram_c3_mode ),
    .dpram_waddr(\m/dram_c3_waddr ),
    .dpram_wclk(\m/dram_c3_wclk ),
    .dpram_we(\m/dram_c3_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c3_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000110),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c3_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c3_di [1:0]),
    .dpram_mode(\m/dram_c3_mode ),
    .dpram_waddr(\m/dram_c3_waddr ),
    .dpram_wclk(\m/dram_c3_wclk ),
    .dpram_we(\m/dram_c3_we ),
    .sr(rst_pad),
    .f(i_data[13:12]),
    .q(\t/busarbitration/instruction [13:12]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c3_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000110),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c3_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c3_di [3:2]),
    .dpram_mode(\m/dram_c3_mode ),
    .dpram_waddr(\m/dram_c3_waddr ),
    .dpram_wclk(\m/dram_c3_wclk ),
    .dpram_we(\m/dram_c3_we ),
    .sr(rst_pad),
    .f(i_data[15:14]),
    .q(\t/busarbitration/instruction [15:14]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c4_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c4_l  (
    .a({o_data[16],n2[0]}),
    .b({o_data[17],n2[1]}),
    .c({o_data[18],n2[2]}),
    .clk(clock_pad),
    .d({o_data[19],n2[3]}),
    .e({open_n19207,memwrite_cs}),
    .dpram_di(\m/dram_c4_di ),
    .dpram_mode(\m/dram_c4_mode ),
    .dpram_waddr(\m/dram_c4_waddr ),
    .dpram_wclk(\m/dram_c4_wclk ),
    .dpram_we(\m/dram_c4_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c4_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c4_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c4_di [1:0]),
    .dpram_mode(\m/dram_c4_mode ),
    .dpram_waddr(\m/dram_c4_waddr ),
    .dpram_wclk(\m/dram_c4_wclk ),
    .dpram_we(\m/dram_c4_we ),
    .sr(rst_pad),
    .f(i_data[17:16]),
    .q(\t/busarbitration/instruction [17:16]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c4_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c4_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c4_di [3:2]),
    .dpram_mode(\m/dram_c4_mode ),
    .dpram_waddr(\m/dram_c4_waddr ),
    .dpram_wclk(\m/dram_c4_wclk ),
    .dpram_we(\m/dram_c4_we ),
    .sr(rst_pad),
    .f(i_data[19:18]),
    .q(\t/busarbitration/instruction [19:18]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c5_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c5_l  (
    .a({o_data[20],n2[0]}),
    .b({o_data[21],n2[1]}),
    .c({o_data[22],n2[2]}),
    .clk(clock_pad),
    .d({o_data[23],n2[3]}),
    .e({open_n19232,memwrite_cs}),
    .dpram_di(\m/dram_c5_di ),
    .dpram_mode(\m/dram_c5_mode ),
    .dpram_waddr(\m/dram_c5_waddr ),
    .dpram_wclk(\m/dram_c5_wclk ),
    .dpram_we(\m/dram_c5_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c5_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c5_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c5_di [1:0]),
    .dpram_mode(\m/dram_c5_mode ),
    .dpram_waddr(\m/dram_c5_waddr ),
    .dpram_wclk(\m/dram_c5_wclk ),
    .dpram_we(\m/dram_c5_we ),
    .sr(rst_pad),
    .f(i_data[21:20]),
    .q(\t/busarbitration/instruction [21:20]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c5_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c5_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c5_di [3:2]),
    .dpram_mode(\m/dram_c5_mode ),
    .dpram_waddr(\m/dram_c5_waddr ),
    .dpram_wclk(\m/dram_c5_wclk ),
    .dpram_we(\m/dram_c5_we ),
    .sr(rst_pad),
    .f(i_data[23:22]),
    .q(\t/busarbitration/instruction [23:22]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c6_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c6_l  (
    .a({o_data[24],n2[0]}),
    .b({o_data[25],n2[1]}),
    .c({o_data[26],n2[2]}),
    .clk(clock_pad),
    .d({o_data[27],n2[3]}),
    .e({open_n19257,memwrite_cs}),
    .dpram_di(\m/dram_c6_di ),
    .dpram_mode(\m/dram_c6_mode ),
    .dpram_waddr(\m/dram_c6_waddr ),
    .dpram_wclk(\m/dram_c6_wclk ),
    .dpram_we(\m/dram_c6_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c6_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c6_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c6_di [1:0]),
    .dpram_mode(\m/dram_c6_mode ),
    .dpram_waddr(\m/dram_c6_waddr ),
    .dpram_wclk(\m/dram_c6_wclk ),
    .dpram_we(\m/dram_c6_we ),
    .sr(rst_pad),
    .f(i_data[25:24]),
    .q(\t/busarbitration/instruction [25:24]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c6_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c6_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c6_di [3:2]),
    .dpram_mode(\m/dram_c6_mode ),
    .dpram_waddr(\m/dram_c6_waddr ),
    .dpram_wclk(\m/dram_c6_wclk ),
    .dpram_we(\m/dram_c6_we ),
    .sr(rst_pad),
    .f(i_data[27:26]),
    .q(\t/busarbitration/instruction [27:26]));
  EG_PHY_LSLICE #(
    //.MACRO("m/dram_c7_l"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \m/dram_c7_l  (
    .a({o_data[28],n2[0]}),
    .b({o_data[29],n2[1]}),
    .c({o_data[30],n2[2]}),
    .clk(clock_pad),
    .d({o_data[31],n2[3]}),
    .e({open_n19282,memwrite_cs}),
    .dpram_di(\m/dram_c7_di ),
    .dpram_mode(\m/dram_c7_mode ),
    .dpram_waddr(\m/dram_c7_waddr ),
    .dpram_wclk(\m/dram_c7_wclk ),
    .dpram_we(\m/dram_c7_we ));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c7_l"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000100),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c7_m0  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c7_di [1:0]),
    .dpram_mode(\m/dram_c7_mode ),
    .dpram_waddr(\m/dram_c7_waddr ),
    .dpram_wclk(\m/dram_c7_wclk ),
    .dpram_we(\m/dram_c7_we ),
    .sr(rst_pad),
    .f(i_data[29:28]),
    .q(\t/busarbitration/instruction [29:28]));
  EG_PHY_MSLICE #(
    //.MACRO("m/dram_c7_l"),
    //.R_POSITION("X0Y0Z1"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000110),
    .INIT_LUT1(16'b0000000000000100),
    .MODE("DPRAM"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMUX("INV"))
    \m/dram_c7_m1  (
    .a({n3[0],n3[0]}),
    .b({n3[1],n3[1]}),
    .c({n3[2],n3[2]}),
    .ce(\t/busarbitration/n3 ),
    .clk(clock_pad),
    .d({n3[3],n3[3]}),
    .dpram_di(\m/dram_c7_di [3:2]),
    .dpram_mode(\m/dram_c7_mode ),
    .dpram_waddr(\m/dram_c7_waddr ),
    .dpram_wclk(\m/dram_c7_wclk ),
    .dpram_we(\m/dram_c7_we ),
    .sr(rst_pad),
    .f(i_data[31:30]),
    .q(\t/busarbitration/instruction [31:30]));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u11_al_u2928  (
    .a({\t/a/EX_A [13],\t/a/EX_A [11]}),
    .b({\t/a/EX_A [14],\t/a/EX_A [12]}),
    .c(2'b00),
    .d({\t/a/EX_B [13],\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/EX_B [14],\t/a/EX_B [12]}),
    .fci(\t/a/alu/add0/c11 ),
    .f({\t/a/alu/n5 [13],\t/a/alu/n5 [11]}),
    .fco(\t/a/alu/add0/c15 ),
    .fx({\t/a/alu/n5 [14],\t/a/alu/n5 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u15_al_u2929  (
    .a({\t/a/EX_A [17],\t/a/EX_A [15]}),
    .b({\t/a/EX_A [18],\t/a/EX_A [16]}),
    .c(2'b00),
    .d({\t/a/EX_B [17],\t/a/EX_B [15]}),
    .e({\t/a/EX_B [18],\t/a/EX_B [16]}),
    .fci(\t/a/alu/add0/c15 ),
    .f({\t/a/alu/n5 [17],\t/a/alu/n5 [15]}),
    .fco(\t/a/alu/add0/c19 ),
    .fx({\t/a/alu/n5 [18],\t/a/alu/n5 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u19_al_u2930  (
    .a({\t/a/EX_A [21],\t/a/EX_A [19]}),
    .b({\t/a/EX_A [22],\t/a/EX_A [20]}),
    .c(2'b00),
    .d({\t/a/EX_B [21],\t/a/EX_B [19]}),
    .e({\t/a/EX_B [22],\t/a/EX_B [20]}),
    .fci(\t/a/alu/add0/c19 ),
    .f({\t/a/alu/n5 [21],\t/a/alu/n5 [19]}),
    .fco(\t/a/alu/add0/c23 ),
    .fx({\t/a/alu/n5 [22],\t/a/alu/n5 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u23_al_u2931  (
    .a({\t/a/EX_A [25],\t/a/EX_A [23]}),
    .b({\t/a/EX_A [26],\t/a/EX_A [24]}),
    .c(2'b00),
    .d({\t/a/EX_B [25],\t/a/EX_B [23]}),
    .e({\t/a/EX_B [26],\t/a/EX_B [24]}),
    .fci(\t/a/alu/add0/c23 ),
    .f({\t/a/alu/n5 [25],\t/a/alu/n5 [23]}),
    .fco(\t/a/alu/add0/c27 ),
    .fx({\t/a/alu/n5 [26],\t/a/alu/n5 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u27_al_u2932  (
    .a({\t/a/EX_A [29],\t/a/EX_A [27]}),
    .b({\t/a/EX_A [30],\t/a/EX_A [28]}),
    .c(2'b00),
    .d({\t/a/EX_B [29],\t/a/EX_B [27]}),
    .e({\t/a/EX_B [30],\t/a/EX_B [28]}),
    .fci(\t/a/alu/add0/c27 ),
    .f({\t/a/alu/n5 [29],\t/a/alu/n5 [27]}),
    .fco(\t/a/alu/add0/c31 ),
    .fx({\t/a/alu/n5 [30],\t/a/alu/n5 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u31_al_u2933  (
    .a({open_n19396,\t/a/EX_A [31]}),
    .c(2'b00),
    .d({open_n19401,\t/a/EX_B [31]}),
    .fci(\t/a/alu/add0/c31 ),
    .f({open_n19418,\t/a/alu/n5 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u3_al_u2926  (
    .a({\t/a/EX_A [5],\t/a/EX_A [3]}),
    .b({\t/a/EX_A [6],\t/a/EX_A [4]}),
    .c(2'b00),
    .d({\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/add0/c3 ),
    .f({\t/a/alu/n5 [5],\t/a/alu/n5 [3]}),
    .fco(\t/a/alu/add0/c7 ),
    .fx({\t/a/alu/n5 [6],\t/a/alu/n5 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/u7_al_u2927  (
    .a({\t/a/EX_A [9],\t/a/EX_A [7]}),
    .b({\t/a/EX_A [10],\t/a/EX_A [8]}),
    .c(2'b00),
    .d({\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/add0/c7 ),
    .f({\t/a/alu/n5 [9],\t/a/alu/n5 [7]}),
    .fco(\t/a/alu/add0/c11 ),
    .fx({\t/a/alu/n5 [10],\t/a/alu/n5 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/add0/ucin_al_u2925"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/add0/ucin_al_u2925  (
    .a({\t/a/EX_A [1],1'b0}),
    .b({\t/a/EX_A [2],\t/a/EX_A [0]}),
    .c(2'b00),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,1'b1}),
    .e({\t/a/EX_B [2],\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({\t/a/alu/n5 [1],open_n19477}),
    .fco(\t/a/alu/add0/c3 ),
    .fx({\t/a/alu/n5 [2],\t/a/alu/n5 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_0|t/a/alu/lt0_cin  (
    .a({\t/a/EX_A [0],1'b0}),
    .b({\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ,open_n19480}),
    .fco(\t/a/alu/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_10|t/a/alu/lt0_9  (
    .a(\t/a/EX_A [10:9]),
    .b({\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/lt0_c9 ),
    .fco(\t/a/alu/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_12|t/a/alu/lt0_11  (
    .a(\t/a/EX_A [12:11]),
    .b({\t/a/EX_B [12],\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/lt0_c11 ),
    .fco(\t/a/alu/lt0_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_14|t/a/alu/lt0_13  (
    .a(\t/a/EX_A [14:13]),
    .b(\t/a/EX_B [14:13]),
    .fci(\t/a/alu/lt0_c13 ),
    .fco(\t/a/alu/lt0_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_16|t/a/alu/lt0_15  (
    .a(\t/a/EX_A [16:15]),
    .b(\t/a/EX_B [16:15]),
    .fci(\t/a/alu/lt0_c15 ),
    .fco(\t/a/alu/lt0_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_18|t/a/alu/lt0_17  (
    .a(\t/a/EX_A [18:17]),
    .b(\t/a/EX_B [18:17]),
    .fci(\t/a/alu/lt0_c17 ),
    .fco(\t/a/alu/lt0_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_20|t/a/alu/lt0_19  (
    .a(\t/a/EX_A [20:19]),
    .b(\t/a/EX_B [20:19]),
    .fci(\t/a/alu/lt0_c19 ),
    .fco(\t/a/alu/lt0_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_22|t/a/alu/lt0_21  (
    .a(\t/a/EX_A [22:21]),
    .b(\t/a/EX_B [22:21]),
    .fci(\t/a/alu/lt0_c21 ),
    .fco(\t/a/alu/lt0_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_24|t/a/alu/lt0_23  (
    .a(\t/a/EX_A [24:23]),
    .b(\t/a/EX_B [24:23]),
    .fci(\t/a/alu/lt0_c23 ),
    .fco(\t/a/alu/lt0_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_26|t/a/alu/lt0_25  (
    .a(\t/a/EX_A [26:25]),
    .b(\t/a/EX_B [26:25]),
    .fci(\t/a/alu/lt0_c25 ),
    .fco(\t/a/alu/lt0_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_28|t/a/alu/lt0_27  (
    .a(\t/a/EX_A [28:27]),
    .b(\t/a/EX_B [28:27]),
    .fci(\t/a/alu/lt0_c27 ),
    .fco(\t/a/alu/lt0_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_2|t/a/alu/lt0_1  (
    .a(\t/a/EX_A [2:1]),
    .b({\t/a/EX_B [2],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/lt0_c1 ),
    .fco(\t/a/alu/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_30|t/a/alu/lt0_29  (
    .a(\t/a/EX_A [30:29]),
    .b(\t/a/EX_B [30:29]),
    .fci(\t/a/alu/lt0_c29 ),
    .fco(\t/a/alu/lt0_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_4|t/a/alu/lt0_3  (
    .a(\t/a/EX_A [4:3]),
    .b({\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/lt0_c3 ),
    .fco(\t/a/alu/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_6|t/a/alu/lt0_5  (
    .a(\t/a/EX_A [6:5]),
    .b({\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/lt0_c5 ),
    .fco(\t/a/alu/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_8|t/a/alu/lt0_7  (
    .a(\t/a/EX_A [8:7]),
    .b({\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/lt0_c7 ),
    .fco(\t/a/alu/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/alu/lt0_0|t/a/alu/lt0_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/alu/lt0_cout|t/a/alu/lt0_31  (
    .a({1'b0,\t/a/EX_A [31]}),
    .b({1'b1,\t/a/EX_B [31]}),
    .fci(\t/a/alu/lt0_c31 ),
    .f({\t/a/alu/n8 ,open_n19884}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u11_al_u2937  (
    .a({\t/a/EX_A [13],\t/a/EX_A [11]}),
    .b({\t/a/EX_A [14],\t/a/EX_A [12]}),
    .c(2'b11),
    .d({\t/a/EX_B [13],\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/EX_B [14],\t/a/EX_B [12]}),
    .fci(\t/a/alu/sub0/c11 ),
    .f({\t/a/alu/n6 [13],\t/a/alu/n6 [11]}),
    .fco(\t/a/alu/sub0/c15 ),
    .fx({\t/a/alu/n6 [14],\t/a/alu/n6 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u15_al_u2938  (
    .a({\t/a/EX_A [17],\t/a/EX_A [15]}),
    .b({\t/a/EX_A [18],\t/a/EX_A [16]}),
    .c(2'b11),
    .d({\t/a/EX_B [17],\t/a/EX_B [15]}),
    .e({\t/a/EX_B [18],\t/a/EX_B [16]}),
    .fci(\t/a/alu/sub0/c15 ),
    .f({\t/a/alu/n6 [17],\t/a/alu/n6 [15]}),
    .fco(\t/a/alu/sub0/c19 ),
    .fx({\t/a/alu/n6 [18],\t/a/alu/n6 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u19_al_u2939  (
    .a({\t/a/EX_A [21],\t/a/EX_A [19]}),
    .b({\t/a/EX_A [22],\t/a/EX_A [20]}),
    .c(2'b11),
    .d({\t/a/EX_B [21],\t/a/EX_B [19]}),
    .e({\t/a/EX_B [22],\t/a/EX_B [20]}),
    .fci(\t/a/alu/sub0/c19 ),
    .f({\t/a/alu/n6 [21],\t/a/alu/n6 [19]}),
    .fco(\t/a/alu/sub0/c23 ),
    .fx({\t/a/alu/n6 [22],\t/a/alu/n6 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u23_al_u2940  (
    .a({\t/a/EX_A [25],\t/a/EX_A [23]}),
    .b({\t/a/EX_A [26],\t/a/EX_A [24]}),
    .c(2'b11),
    .d({\t/a/EX_B [25],\t/a/EX_B [23]}),
    .e({\t/a/EX_B [26],\t/a/EX_B [24]}),
    .fci(\t/a/alu/sub0/c23 ),
    .f({\t/a/alu/n6 [25],\t/a/alu/n6 [23]}),
    .fco(\t/a/alu/sub0/c27 ),
    .fx({\t/a/alu/n6 [26],\t/a/alu/n6 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u27_al_u2941  (
    .a({\t/a/EX_A [29],\t/a/EX_A [27]}),
    .b({\t/a/EX_A [30],\t/a/EX_A [28]}),
    .c(2'b11),
    .d({\t/a/EX_B [29],\t/a/EX_B [27]}),
    .e({\t/a/EX_B [30],\t/a/EX_B [28]}),
    .fci(\t/a/alu/sub0/c27 ),
    .f({\t/a/alu/n6 [29],\t/a/alu/n6 [27]}),
    .fco(\t/a/alu/sub0/c31 ),
    .fx({\t/a/alu/n6 [30],\t/a/alu/n6 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u31_al_u2942  (
    .a({open_n19980,\t/a/EX_A [31]}),
    .c(2'b11),
    .d({open_n19985,\t/a/EX_B [31]}),
    .fci(\t/a/alu/sub0/c31 ),
    .f({open_n20002,\t/a/alu/n6 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u3_al_u2935  (
    .a({\t/a/EX_A [5],\t/a/EX_A [3]}),
    .b({\t/a/EX_A [6],\t/a/EX_A [4]}),
    .c(2'b11),
    .d({\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/sub0/c3 ),
    .f({\t/a/alu/n6 [5],\t/a/alu/n6 [3]}),
    .fco(\t/a/alu/sub0/c7 ),
    .fx({\t/a/alu/n6 [6],\t/a/alu/n6 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/u7_al_u2936  (
    .a({\t/a/EX_A [9],\t/a/EX_A [7]}),
    .b({\t/a/EX_A [10],\t/a/EX_A [8]}),
    .c(2'b11),
    .d({\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o }),
    .e({\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o }),
    .fci(\t/a/alu/sub0/c7 ),
    .f({\t/a/alu/n6 [9],\t/a/alu/n6 [7]}),
    .fco(\t/a/alu/sub0/c11 ),
    .fx({\t/a/alu/n6 [10],\t/a/alu/n6 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/alu/sub0/ucin_al_u2934"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/alu/sub0/ucin_al_u2934  (
    .a({\t/a/EX_A [1],1'b0}),
    .b({\t/a/EX_A [2],\t/a/EX_A [0]}),
    .c(2'b11),
    .d({\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,1'b1}),
    .e({\t/a/EX_B [2],\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .f({\t/a/alu/n6 [1],open_n20061}),
    .fco(\t/a/alu/sub0/c3 ),
    .fx({\t/a/alu/n6 [2],\t/a/alu/n6 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u11_al_u2946  (
    .a({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .b({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [13],\t/a/ID_jump_regdat1 [11]}),
    .e({\t/a/ID_jump_regdat1 [14],\t/a/ID_jump_regdat1 [12]}),
    .fci(\t/a/condition/add0/c11 ),
    .f({\t/a/condition/n5 [13],\t/a/condition/n5 [11]}),
    .fco(\t/a/condition/add0/c15 ),
    .fx({\t/a/condition/n5 [14],\t/a/condition/n5 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u15_al_u2947  (
    .a({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .b({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [17],\t/a/ID_jump_regdat1 [15]}),
    .e({\t/a/ID_jump_regdat1 [18],\t/a/ID_jump_regdat1 [16]}),
    .fci(\t/a/condition/add0/c15 ),
    .f({\t/a/condition/n5 [17],\t/a/condition/n5 [15]}),
    .fco(\t/a/condition/add0/c19 ),
    .fx({\t/a/condition/n5 [18],\t/a/condition/n5 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u19_al_u2948  (
    .a({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .b({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [21],\t/a/ID_jump_regdat1 [19]}),
    .e({\t/a/ID_jump_regdat1 [22],\t/a/ID_jump_regdat1 [20]}),
    .fci(\t/a/condition/add0/c19 ),
    .f({\t/a/condition/n5 [21],\t/a/condition/n5 [19]}),
    .fco(\t/a/condition/add0/c23 ),
    .fx({\t/a/condition/n5 [22],\t/a/condition/n5 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u23_al_u2949  (
    .a({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .b({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [25],\t/a/ID_jump_regdat1 [23]}),
    .e({\t/a/ID_jump_regdat1 [26],\t/a/ID_jump_regdat1 [24]}),
    .fci(\t/a/condition/add0/c23 ),
    .f({\t/a/condition/n5 [25],\t/a/condition/n5 [23]}),
    .fco(\t/a/condition/add0/c27 ),
    .fx({\t/a/condition/n5 [26],\t/a/condition/n5 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u27_al_u2950  (
    .a({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .b({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [29],\t/a/ID_jump_regdat1 [27]}),
    .e({\t/a/ID_jump_regdat1 [30],\t/a/ID_jump_regdat1 [28]}),
    .fci(\t/a/condition/add0/c27 ),
    .f({\t/a/condition/n5 [29],\t/a/condition/n5 [27]}),
    .fco(\t/a/condition/add0/c31 ),
    .fx({\t/a/condition/n5 [30],\t/a/condition/n5 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u31_al_u2951  (
    .a({open_n20154,\t/a/ID_fun7 [6]}),
    .c(2'b00),
    .d({open_n20159,\t/a/ID_jump_regdat1 [31]}),
    .fci(\t/a/condition/add0/c31 ),
    .f({open_n20176,\t/a/condition/n5 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u3_al_u2944  (
    .a({\t/a/ID_fun7 [0],\t/a/ID_rs2 [3]}),
    .b({\t/a/ID_fun7 [1],\t/a/ID_rs2 [4]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [5],\t/a/ID_jump_regdat1 [3]}),
    .e({\t/a/ID_jump_regdat1 [6],\t/a/ID_jump_regdat1 [4]}),
    .fci(\t/a/condition/add0/c3 ),
    .f({\t/a/condition/n5 [5],\t/a/condition/n5 [3]}),
    .fco(\t/a/condition/add0/c7 ),
    .fx({\t/a/condition/n5 [6],\t/a/condition/n5 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/u7_al_u2945  (
    .a({\t/a/ID_fun7 [4],\t/a/ID_fun7 [2]}),
    .b({\t/a/ID_fun7 [5],\t/a/ID_fun7 [3]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [9],\t/a/ID_jump_regdat1 [7]}),
    .e({\t/a/ID_jump_regdat1 [10],\t/a/ID_jump_regdat1 [8]}),
    .fci(\t/a/condition/add0/c7 ),
    .f({\t/a/condition/n5 [9],\t/a/condition/n5 [7]}),
    .fco(\t/a/condition/add0/c11 ),
    .fx({\t/a/condition/n5 [10],\t/a/condition/n5 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/condition/add0/ucin_al_u2943"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/condition/add0/ucin_al_u2943  (
    .a({\t/a/ID_rs2 [1],1'b0}),
    .b({\t/a/ID_rs2 [2],\t/a/ID_rs2 [0]}),
    .c(2'b00),
    .d({\t/a/ID_jump_regdat1 [1],1'b1}),
    .e({\t/a/ID_jump_regdat1 [2],\t/a/ID_jump_regdat1 [0]}),
    .f({\t/a/condition/n5 [1],open_n20235}),
    .fco(\t/a/condition/add0/c3 ),
    .fx({\t/a/condition/n5 [2],open_n20236}));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_0|t/a/condition/lt0_cin  (
    .a({\t/a/ID_jump_regdat1 [0],1'b0}),
    .b({\t/a/ID_jump_regdat2 [0],open_n20239}),
    .fco(\t/a/condition/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_10|t/a/condition/lt0_9  (
    .a(\t/a/ID_jump_regdat1 [10:9]),
    .b(\t/a/ID_jump_regdat2 [10:9]),
    .fci(\t/a/condition/lt0_c9 ),
    .fco(\t/a/condition/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_12|t/a/condition/lt0_11  (
    .a(\t/a/ID_jump_regdat1 [12:11]),
    .b(\t/a/ID_jump_regdat2 [12:11]),
    .fci(\t/a/condition/lt0_c11 ),
    .fco(\t/a/condition/lt0_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_14|t/a/condition/lt0_13  (
    .a(\t/a/ID_jump_regdat1 [14:13]),
    .b(\t/a/ID_jump_regdat2 [14:13]),
    .fci(\t/a/condition/lt0_c13 ),
    .fco(\t/a/condition/lt0_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_16|t/a/condition/lt0_15  (
    .a(\t/a/ID_jump_regdat1 [16:15]),
    .b(\t/a/ID_jump_regdat2 [16:15]),
    .fci(\t/a/condition/lt0_c15 ),
    .fco(\t/a/condition/lt0_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_18|t/a/condition/lt0_17  (
    .a(\t/a/ID_jump_regdat1 [18:17]),
    .b(\t/a/ID_jump_regdat2 [18:17]),
    .fci(\t/a/condition/lt0_c17 ),
    .fco(\t/a/condition/lt0_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_20|t/a/condition/lt0_19  (
    .a(\t/a/ID_jump_regdat1 [20:19]),
    .b(\t/a/ID_jump_regdat2 [20:19]),
    .fci(\t/a/condition/lt0_c19 ),
    .fco(\t/a/condition/lt0_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_22|t/a/condition/lt0_21  (
    .a(\t/a/ID_jump_regdat1 [22:21]),
    .b(\t/a/ID_jump_regdat2 [22:21]),
    .fci(\t/a/condition/lt0_c21 ),
    .fco(\t/a/condition/lt0_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_24|t/a/condition/lt0_23  (
    .a(\t/a/ID_jump_regdat1 [24:23]),
    .b(\t/a/ID_jump_regdat2 [24:23]),
    .fci(\t/a/condition/lt0_c23 ),
    .fco(\t/a/condition/lt0_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_26|t/a/condition/lt0_25  (
    .a(\t/a/ID_jump_regdat1 [26:25]),
    .b(\t/a/ID_jump_regdat2 [26:25]),
    .fci(\t/a/condition/lt0_c25 ),
    .fco(\t/a/condition/lt0_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_28|t/a/condition/lt0_27  (
    .a(\t/a/ID_jump_regdat1 [28:27]),
    .b(\t/a/ID_jump_regdat2 [28:27]),
    .fci(\t/a/condition/lt0_c27 ),
    .fco(\t/a/condition/lt0_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_2|t/a/condition/lt0_1  (
    .a(\t/a/ID_jump_regdat1 [2:1]),
    .b(\t/a/ID_jump_regdat2 [2:1]),
    .fci(\t/a/condition/lt0_c1 ),
    .fco(\t/a/condition/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_30|t/a/condition/lt0_29  (
    .a(\t/a/ID_jump_regdat1 [30:29]),
    .b(\t/a/ID_jump_regdat2 [30:29]),
    .fci(\t/a/condition/lt0_c29 ),
    .fco(\t/a/condition/lt0_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_4|t/a/condition/lt0_3  (
    .a(\t/a/ID_jump_regdat1 [4:3]),
    .b(\t/a/ID_jump_regdat2 [4:3]),
    .fci(\t/a/condition/lt0_c3 ),
    .fco(\t/a/condition/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_6|t/a/condition/lt0_5  (
    .a(\t/a/ID_jump_regdat1 [6:5]),
    .b(\t/a/ID_jump_regdat2 [6:5]),
    .fci(\t/a/condition/lt0_c5 ),
    .fco(\t/a/condition/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_8|t/a/condition/lt0_7  (
    .a(\t/a/ID_jump_regdat1 [8:7]),
    .b(\t/a/ID_jump_regdat2 [8:7]),
    .fci(\t/a/condition/lt0_c7 ),
    .fco(\t/a/condition/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt0_0|t/a/condition/lt0_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt0_cout|t/a/condition/lt0_31  (
    .a({1'b0,\t/a/ID_jump_regdat1 [31]}),
    .b({1'b1,\t/a/ID_jump_regdat2 [31]}),
    .fci(\t/a/condition/lt0_c31 ),
    .f({\t/a/condition/n9 ,open_n20643}));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_0|t/a/condition/lt1_cin  (
    .a({\t/a/ID_jump_regdat1 [0],1'b0}),
    .b({\t/a/ID_jump_regdat2 [0],open_n20649}),
    .fco(\t/a/condition/lt1_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_10|t/a/condition/lt1_9  (
    .a(\t/a/ID_jump_regdat1 [10:9]),
    .b(\t/a/ID_jump_regdat2 [10:9]),
    .fci(\t/a/condition/lt1_c9 ),
    .fco(\t/a/condition/lt1_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_12|t/a/condition/lt1_11  (
    .a(\t/a/ID_jump_regdat1 [12:11]),
    .b(\t/a/ID_jump_regdat2 [12:11]),
    .fci(\t/a/condition/lt1_c11 ),
    .fco(\t/a/condition/lt1_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_14|t/a/condition/lt1_13  (
    .a(\t/a/ID_jump_regdat1 [14:13]),
    .b(\t/a/ID_jump_regdat2 [14:13]),
    .fci(\t/a/condition/lt1_c13 ),
    .fco(\t/a/condition/lt1_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_16|t/a/condition/lt1_15  (
    .a(\t/a/ID_jump_regdat1 [16:15]),
    .b(\t/a/ID_jump_regdat2 [16:15]),
    .fci(\t/a/condition/lt1_c15 ),
    .fco(\t/a/condition/lt1_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_18|t/a/condition/lt1_17  (
    .a(\t/a/ID_jump_regdat1 [18:17]),
    .b(\t/a/ID_jump_regdat2 [18:17]),
    .fci(\t/a/condition/lt1_c17 ),
    .fco(\t/a/condition/lt1_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_20|t/a/condition/lt1_19  (
    .a(\t/a/ID_jump_regdat1 [20:19]),
    .b(\t/a/ID_jump_regdat2 [20:19]),
    .fci(\t/a/condition/lt1_c19 ),
    .fco(\t/a/condition/lt1_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_22|t/a/condition/lt1_21  (
    .a(\t/a/ID_jump_regdat1 [22:21]),
    .b(\t/a/ID_jump_regdat2 [22:21]),
    .fci(\t/a/condition/lt1_c21 ),
    .fco(\t/a/condition/lt1_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_24|t/a/condition/lt1_23  (
    .a(\t/a/ID_jump_regdat1 [24:23]),
    .b(\t/a/ID_jump_regdat2 [24:23]),
    .fci(\t/a/condition/lt1_c23 ),
    .fco(\t/a/condition/lt1_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_26|t/a/condition/lt1_25  (
    .a(\t/a/ID_jump_regdat1 [26:25]),
    .b(\t/a/ID_jump_regdat2 [26:25]),
    .fci(\t/a/condition/lt1_c25 ),
    .fco(\t/a/condition/lt1_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_28|t/a/condition/lt1_27  (
    .a(\t/a/ID_jump_regdat1 [28:27]),
    .b(\t/a/ID_jump_regdat2 [28:27]),
    .fci(\t/a/condition/lt1_c27 ),
    .fco(\t/a/condition/lt1_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_2|t/a/condition/lt1_1  (
    .a(\t/a/ID_jump_regdat1 [2:1]),
    .b(\t/a/ID_jump_regdat2 [2:1]),
    .fci(\t/a/condition/lt1_c1 ),
    .fco(\t/a/condition/lt1_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_30|t/a/condition/lt1_29  (
    .a(\t/a/ID_jump_regdat1 [30:29]),
    .b(\t/a/ID_jump_regdat2 [30:29]),
    .fci(\t/a/condition/lt1_c29 ),
    .fco(\t/a/condition/lt1_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_4|t/a/condition/lt1_3  (
    .a(\t/a/ID_jump_regdat1 [4:3]),
    .b(\t/a/ID_jump_regdat2 [4:3]),
    .fci(\t/a/condition/lt1_c3 ),
    .fco(\t/a/condition/lt1_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_6|t/a/condition/lt1_5  (
    .a(\t/a/ID_jump_regdat1 [6:5]),
    .b(\t/a/ID_jump_regdat2 [6:5]),
    .fci(\t/a/condition/lt1_c5 ),
    .fco(\t/a/condition/lt1_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_8|t/a/condition/lt1_7  (
    .a(\t/a/ID_jump_regdat1 [8:7]),
    .b(\t/a/ID_jump_regdat2 [8:7]),
    .fci(\t/a/condition/lt1_c7 ),
    .fco(\t/a/condition/lt1_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("t/a/condition/lt1_0|t/a/condition/lt1_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \t/a/condition/lt1_cout_al_u2977  (
    .a({open_n21035,1'b0}),
    .b({open_n21036,1'b1}),
    .fci(\t/a/condition/lt1_c31 ),
    .f({open_n21055,\t/a/condition/n10 }));
  // flow_line_reg.v(234)
  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg0_b1|t/a/mem_wb/reg2_b1  (
    .a({\t/a/aluin/n12_lutinv ,\t/a/MEM_rd [1]}),
    .b({_al_u1984_o,\t/a/MEM_rd [4]}),
    .c({\t/a/EX_rs2 [1],\t/a/EX_rs2 [1]}),
    .clk(clock_pad),
    .d({\t/a/EX_rd [1],\t/a/EX_rs2 [4]}),
    .mi({\t/a/EX_rd [1],\t/a/MEM_rd [1]}),
    .sr(rst_pad),
    .f({_al_u2073_o,_al_u1969_o}),
    .q({\t/a/MEM_rd [1],\t/a/WB_rd [1]}));  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(~C*A))"),
    //.LUTF1("(~(C*B)*~(D*A))"),
    //.LUTG0("(~(D*~B)*~(~C*A))"),
    //.LUTG1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100010011110101),
    .INIT_LUTF1(16'b0001010100111111),
    .INIT_LUTG0(16'b1100010011110101),
    .INIT_LUTG1(16'b0001010100111111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg0_b3|t/a/mem_wb/reg2_b3  (
    .a({\t/a/aluin/n12_lutinv ,\t/a/MEM_rd [3]}),
    .b({_al_u1984_o,\t/a/MEM_rd [4]}),
    .c({\t/a/EX_rs2 [3],\t/a/EX_rs2 [3]}),
    .clk(clock_pad),
    .d({\t/a/EX_rd [3],\t/a/EX_rs2 [4]}),
    .mi({\t/a/EX_rd [3],\t/a/MEM_rd [3]}),
    .sr(rst_pad),
    .f({_al_u2010_o,_al_u1970_o}),
    .q({\t/a/MEM_rd [3],\t/a/WB_rd [3]}));  // flow_line_reg.v(234)
  // flow_line_reg.v(139)
  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*C))"),
    //.LUT1("(~(C*B)*~(D*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111011101110),
    .INIT_LUT1(16'b0001010100111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg0_b4|t/a/id_ex/reg3_b4  (
    .a({\t/a/aluin/n12_lutinv ,\t/a/aluin/sel1_b24/B9 }),
    .b({_al_u1984_o,_al_u2007_o}),
    .c({\t/a/EX_rs2 [4],_al_u1803_o}),
    .clk(clock_pad),
    .d({\t/a/EX_rd [4],\t/a/EX_rs2 [4]}),
    .mi({\t/a/EX_rd [4],\t/a/ID_rs2 [4]}),
    .sr(rst_pad),
    .f({_al_u2000_o,\t/a/EX_B [24]}),
    .q({\t/a/MEM_rd [4],\t/a/EX_rs2 [4]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b0011001100001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg1_b2|t/a/id_ex/reg0_b2  (
    .a({open_n21111,_al_u1049_o}),
    .b({\t/a/MEM_aludat [2],_al_u1248_o}),
    .c({\t/a/EX_regdat2 [2],_al_u1258_o}),
    .clk(clock_pad),
    .d({\t/a/alu_B_select [0],\t/a/reg_writedat [2]}),
    .mi({\t/a/EX_regdat2 [2],open_n21123}),
    .sr(rst_pad),
    .f({_al_u2092_o,\t/a/ID_read_dat2 [2]}),
    .q({\t/a/MEM_regdat2 [2],\t/a/EX_regdat2 [2]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(~C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg2_b1|t/a/id_ex/reg6_b1  (
    .a({open_n21127,_al_u1747_o}),
    .b({\t/a/EX_op [1],\t/a/ID_op [0]}),
    .c({\t/a/EX_op [2],\t/a/ID_op [1]}),
    .clk(clock_pad),
    .d({\t/a/EX_op [0],\t/a/ID_op [2]}),
    .mi({\t/a/EX_op [1],\t/a/ID_op [1]}),
    .sr(rst_pad),
    .f({_al_u1739_o,\t/a/condition/sel1/B2 }),
    .q({\t/a/MEM_op [1],\t/a/EX_op [1]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg2_b2|t/a/ex_mem/reg2_b0  (
    .b({\t/a/MEM_op [1],\t/a/EX_op [1]}),
    .c({\t/a/MEM_op [2],\t/a/EX_op [2]}),
    .clk(clock_pad),
    .d({\t/a/MEM_op [0],\t/a/EX_op [0]}),
    .mi({\t/a/EX_op [2],\t/a/EX_op [0]}),
    .sr(rst_pad),
    .f({_al_u290_o,_al_u1801_o}),
    .q({\t/a/MEM_op [2],\t/a/MEM_op [0]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*D*C*~B*A)"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("(~1*D*C*~B*A)"),
    //.LUTG1("(~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000000000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg2_b3|t/a/id_ex/reg6_b6  (
    .a({_al_u1739_o,_al_u1739_o}),
    .b({\t/a/EX_op [3],\t/a/EX_op [3]}),
    .c(\t/a/EX_op [5:4]),
    .clk(clock_pad),
    .d(\t/a/EX_op [6:5]),
    .e({open_n21163,\t/a/EX_op [6]}),
    .mi({\t/a/EX_op [3],\t/a/ID_op [6]}),
    .sr(rst_pad),
    .f({_al_u1984_o,\t/a/aluin/n10_lutinv }),
    .q({\t/a/MEM_op [3],\t/a/EX_op [6]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(191)
  EG_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*B*A)"),
    //.LUTF1("(C*~(~B*~(D*A)))"),
    //.LUTG0("(~1*~D*~C*B*A)"),
    //.LUTG1("(C*~(~B*~(D*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b1110000011000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1110000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg3_b2|t/a/id_ex/reg1_b2  (
    .a({_al_u1984_o,\t/a/aluin/n35_lutinv }),
    .b({\t/a/aluin/n10_lutinv ,\t/a/aluin/n10_lutinv }),
    .c({\t/a/EX_fun3 [2],\t/a/EX_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/EX_op [4],\t/a/EX_fun3 [1]}),
    .e({open_n21180,\t/a/EX_fun3 [2]}),
    .mi({\t/a/EX_fun3 [2],\t/a/ID_fun3 [2]}),
    .sr(rst_pad),
    .f({\t/a/EX_operation [2],_al_u2126_o}),
    .q({\t/a/MEM_fun3 [2],\t/a/EX_fun3 [2]}));  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(~C*~(~D*~A))))"),
    //.LUT1("(B*~(1*~(~C*~(~D*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000110000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b1  (
    .a({\t/a/alu/mux0_b1/B1_0 ,\t/a/alu/mux0_b1/B1_0 }),
    .b({_al_u2586_o,_al_u2586_o}),
    .c({_al_u2587_o,_al_u2587_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n21207,_al_u2128_o}),
    .sr(rst_pad),
    .fx({open_n21211,\t/a/aludat [1]}),
    .q({open_n21212,\t/a/MEM_aludat [1]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b10  (
    .a({_al_u2478_o,_al_u2478_o}),
    .b({_al_u2480_o,_al_u2480_o}),
    .c({_al_u2486_o,_al_u2486_o}),
    .clk(clock_pad),
    .d({_al_u2279_o,_al_u2279_o}),
    .mi({open_n21224,_al_u2161_o}),
    .sr(rst_pad),
    .q({open_n21230,\t/a/MEM_aludat [10]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b11  (
    .a({_al_u2468_o,_al_u2468_o}),
    .b({_al_u2470_o,_al_u2470_o}),
    .c({_al_u2476_o,_al_u2476_o}),
    .clk(clock_pad),
    .d({_al_u2262_o,_al_u2262_o}),
    .mi({open_n21242,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n21246,\t/a/aludat [11]}),
    .q({open_n21247,\t/a/MEM_aludat [11]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b12  (
    .a({_al_u2458_o,_al_u2458_o}),
    .b({_al_u2460_o,_al_u2460_o}),
    .c({_al_u2466_o,_al_u2466_o}),
    .clk(clock_pad),
    .d({_al_u2242_o,_al_u2242_o}),
    .mi({open_n21259,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n21263,\t/a/aludat [12]}),
    .q({open_n21264,\t/a/MEM_aludat [12]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b13  (
    .a({_al_u2448_o,_al_u2448_o}),
    .b({_al_u2450_o,_al_u2450_o}),
    .c({_al_u2456_o,_al_u2456_o}),
    .clk(clock_pad),
    .d({_al_u2219_o,_al_u2219_o}),
    .mi({open_n21276,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n21280,\t/a/aludat [13]}),
    .q({open_n21281,\t/a/MEM_aludat [13]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b14  (
    .a({_al_u2438_o,_al_u2438_o}),
    .b({_al_u2440_o,_al_u2440_o}),
    .c({_al_u2446_o,_al_u2446_o}),
    .clk(clock_pad),
    .d({_al_u2187_o,_al_u2187_o}),
    .mi({open_n21293,_al_u2161_o}),
    .sr(rst_pad),
    .q({open_n21299,\t/a/MEM_aludat [14]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b17  (
    .a({_al_u2405_o,_al_u2405_o}),
    .b({_al_u2406_o,_al_u2406_o}),
    .c({_al_u2412_o,_al_u2412_o}),
    .clk(clock_pad),
    .d({_al_u2413_o,_al_u2413_o}),
    .mi({open_n21311,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21315,\t/a/aludat [17]}),
    .q({open_n21316,\t/a/MEM_aludat [17]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~(0*~A))))"),
    //.LUT1("~(~D*~(C*~(B*~(1*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1111111101110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b18  (
    .a({_al_u2392_o,_al_u2392_o}),
    .b({_al_u2393_o,_al_u2393_o}),
    .c({_al_u2399_o,_al_u2399_o}),
    .clk(clock_pad),
    .d({_al_u2400_o,_al_u2400_o}),
    .mi({open_n21328,_al_u2128_o}),
    .sr(rst_pad),
    .fx({open_n21332,\t/a/aludat [18]}),
    .q({open_n21333,\t/a/MEM_aludat [18]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(B*~(0*~A))))"),
    //.LUT1("~(~D*~(C*~(B*~(1*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100110000),
    .INIT_LUT1(16'b1111111101110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b19  (
    .a({_al_u2380_o,_al_u2380_o}),
    .b({_al_u2381_o,_al_u2381_o}),
    .c({_al_u2387_o,_al_u2387_o}),
    .clk(clock_pad),
    .d({_al_u2388_o,_al_u2388_o}),
    .mi({open_n21345,_al_u2128_o}),
    .sr(rst_pad),
    .fx({open_n21349,\t/a/aludat [19]}),
    .q({open_n21350,\t/a/MEM_aludat [19]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(~C*~(~D*~A))))"),
    //.LUT1("(B*~(1*~(~C*~(~D*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000110000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b2  (
    .a({\t/a/alu/mux0_b2/B1_0 ,\t/a/alu/mux0_b2/B1_0 }),
    .b({_al_u2564_o,_al_u2564_o}),
    .c({_al_u2565_o,_al_u2565_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n21362,_al_u2128_o}),
    .sr(rst_pad),
    .fx({open_n21366,\t/a/aludat [2]}),
    .q({open_n21367,\t/a/MEM_aludat [2]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b20  (
    .a({_al_u2368_o,_al_u2368_o}),
    .b({_al_u2369_o,_al_u2369_o}),
    .c({_al_u2375_o,_al_u2375_o}),
    .clk(clock_pad),
    .d({_al_u2376_o,_al_u2376_o}),
    .mi({open_n21379,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21383,\t/a/aludat [20]}),
    .q({open_n21384,\t/a/MEM_aludat [20]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b21  (
    .a({_al_u2355_o,_al_u2355_o}),
    .b({_al_u2356_o,_al_u2356_o}),
    .c({_al_u2362_o,_al_u2362_o}),
    .clk(clock_pad),
    .d({_al_u2363_o,_al_u2363_o}),
    .mi({open_n21396,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21400,\t/a/aludat [21]}),
    .q({open_n21401,\t/a/MEM_aludat [21]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b22  (
    .a({_al_u2342_o,_al_u2342_o}),
    .b({_al_u2343_o,_al_u2343_o}),
    .c({_al_u2349_o,_al_u2349_o}),
    .clk(clock_pad),
    .d({_al_u2350_o,_al_u2350_o}),
    .mi({open_n21413,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21417,\t/a/aludat [22]}),
    .q({open_n21418,\t/a/MEM_aludat [22]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b23  (
    .a({_al_u2329_o,_al_u2329_o}),
    .b({_al_u2330_o,_al_u2330_o}),
    .c({_al_u2336_o,_al_u2336_o}),
    .clk(clock_pad),
    .d({_al_u2337_o,_al_u2337_o}),
    .mi({open_n21430,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21434,\t/a/aludat [23]}),
    .q({open_n21435,\t/a/MEM_aludat [23]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b24  (
    .a({_al_u2310_o,_al_u2310_o}),
    .b({_al_u2317_o,_al_u2317_o}),
    .c({_al_u2323_o,_al_u2323_o}),
    .clk(clock_pad),
    .d({_al_u2324_o,_al_u2324_o}),
    .mi({open_n21447,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21451,\t/a/aludat [24]}),
    .q({open_n21452,\t/a/MEM_aludat [24]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b25  (
    .a({_al_u2293_o,_al_u2293_o}),
    .b({_al_u2301_o,_al_u2301_o}),
    .c({_al_u2307_o,_al_u2307_o}),
    .clk(clock_pad),
    .d({_al_u2308_o,_al_u2308_o}),
    .mi({open_n21464,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21468,\t/a/aludat [25]}),
    .q({open_n21469,\t/a/MEM_aludat [25]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b26  (
    .a({_al_u2276_o,_al_u2276_o}),
    .b({_al_u2284_o,_al_u2284_o}),
    .c({_al_u2290_o,_al_u2290_o}),
    .clk(clock_pad),
    .d({_al_u2291_o,_al_u2291_o}),
    .mi({open_n21481,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21485,\t/a/aludat [26]}),
    .q({open_n21486,\t/a/MEM_aludat [26]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b27  (
    .a({_al_u2259_o,_al_u2259_o}),
    .b({_al_u2267_o,_al_u2267_o}),
    .c({_al_u2273_o,_al_u2273_o}),
    .clk(clock_pad),
    .d({_al_u2274_o,_al_u2274_o}),
    .mi({open_n21498,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21502,\t/a/aludat [27]}),
    .q({open_n21503,\t/a/MEM_aludat [27]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b28  (
    .a({_al_u2236_o,_al_u2236_o}),
    .b({_al_u2250_o,_al_u2250_o}),
    .c({_al_u2256_o,_al_u2256_o}),
    .clk(clock_pad),
    .d({_al_u2257_o,_al_u2257_o}),
    .mi({open_n21515,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21519,\t/a/aludat [28]}),
    .q({open_n21520,\t/a/MEM_aludat [28]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b29  (
    .a({_al_u2212_o,_al_u2212_o}),
    .b({_al_u2227_o,_al_u2227_o}),
    .c({_al_u2233_o,_al_u2233_o}),
    .clk(clock_pad),
    .d({_al_u2234_o,_al_u2234_o}),
    .mi({open_n21532,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21536,\t/a/aludat [29]}),
    .q({open_n21537,\t/a/MEM_aludat [29]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(~C*~(~D*~A))))"),
    //.LUT1("(B*~(1*~(~C*~(~D*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000110000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b3  (
    .a({\t/a/alu/mux0_b3/B1_0 ,\t/a/alu/mux0_b3/B1_0 }),
    .b({_al_u2555_o,_al_u2555_o}),
    .c({_al_u2556_o,_al_u2556_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n21549,_al_u2128_o}),
    .sr(rst_pad),
    .q({open_n21555,\t/a/MEM_aludat [3]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b30  (
    .a({_al_u2172_o,_al_u2172_o}),
    .b({_al_u2203_o,_al_u2203_o}),
    .c({_al_u2209_o,_al_u2209_o}),
    .clk(clock_pad),
    .d({_al_u2210_o,_al_u2210_o}),
    .mi({open_n21567,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21571,\t/a/aludat [30]}),
    .q({open_n21572,\t/a/MEM_aludat [30]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("~(~D*~(C*~(~0*~(~B*~A))))"),
    //.LUT1("~(~D*~(C*~(~1*~(~B*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111100010000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b31  (
    .a({_al_u2130_o,_al_u2130_o}),
    .b({_al_u2163_o,_al_u2163_o}),
    .c({_al_u2168_o,_al_u2168_o}),
    .clk(clock_pad),
    .d({_al_u2170_o,_al_u2170_o}),
    .mi({open_n21584,\t/a/EX_operation [2]}),
    .sr(rst_pad),
    .fx({open_n21588,\t/a/aludat [31]}),
    .q({open_n21589,\t/a/MEM_aludat [31]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(~C*~(~D*~A))))"),
    //.LUT1("(B*~(1*~(~C*~(~D*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000110000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b5  (
    .a({\t/a/alu/mux0_b5/B1_0 ,\t/a/alu/mux0_b5/B1_0 }),
    .b({_al_u2535_o,_al_u2535_o}),
    .c({_al_u2536_o,_al_u2536_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n21601,_al_u2128_o}),
    .sr(rst_pad),
    .q({open_n21607,\t/a/MEM_aludat [5]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(0*~(~C*~(~D*~A))))"),
    //.LUT1("(B*~(1*~(~C*~(~D*~A))))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100110011001100),
    .INIT_LUT1(16'b0000110000001000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b6  (
    .a({\t/a/alu/mux0_b6/B1_0 ,\t/a/alu/mux0_b6/B1_0 }),
    .b({_al_u2525_o,_al_u2525_o}),
    .c({_al_u2526_o,_al_u2526_o}),
    .clk(clock_pad),
    .d({\t/a/EX_operation [2],\t/a/EX_operation [2]}),
    .mi({open_n21619,_al_u2128_o}),
    .sr(rst_pad),
    .q({open_n21625,\t/a/MEM_aludat [6]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*D)))"),
    //.LUT1("(~C*B*~(A*~(1*D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000110000000100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b7  (
    .a({_al_u2508_o,_al_u2508_o}),
    .b({_al_u2510_o,_al_u2510_o}),
    .c({_al_u2516_o,_al_u2516_o}),
    .clk(clock_pad),
    .d({\t/a/alu/n260_lutinv ,\t/a/alu/n260_lutinv }),
    .mi({open_n21637,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n21641,\t/a/aludat [7]}),
    .q({open_n21642,\t/a/MEM_aludat [7]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b8  (
    .a({_al_u2498_o,_al_u2498_o}),
    .b({_al_u2500_o,_al_u2500_o}),
    .c({_al_u2506_o,_al_u2506_o}),
    .clk(clock_pad),
    .d({_al_u2312_o,_al_u2312_o}),
    .mi({open_n21654,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n21658,\t/a/aludat [8]}),
    .q({open_n21659,\t/a/MEM_aludat [8]}));  // flow_line_reg.v(191)
  EG_PHY_MSLICE #(
    //.LUT0("(~C*B*~(A*~(0*~D)))"),
    //.LUT1("(~C*B*~(A*~(1*~D)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010000000100),
    .INIT_LUT1(16'b0000010000001100),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/ex_mem/reg4_b9  (
    .a({_al_u2488_o,_al_u2488_o}),
    .b({_al_u2490_o,_al_u2490_o}),
    .c({_al_u2496_o,_al_u2496_o}),
    .clk(clock_pad),
    .d({_al_u2296_o,_al_u2296_o}),
    .mi({open_n21671,_al_u2161_o}),
    .sr(rst_pad),
    .fx({open_n21675,\t/a/aludat [9]}),
    .q({open_n21676,\t/a/MEM_aludat [9]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b0|t/a/ex_mem/reg1_b0  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1710_o,\t/a/alu_B_select [1]}),
    .c({_al_u1720_o,\t/a/MEM_aludat [0]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [0],\t/a/EX_regdat2 [0]}),
    .mi({open_n21681,\t/a/EX_regdat2 [0]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [0],_al_u2075_o}),
    .q({\t/a/EX_regdat2 [0],\t/a/MEM_regdat2 [0]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b10|t/a/ex_mem/reg1_b10  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1689_o,\t/a/alu_B_select [1]}),
    .c({_al_u1699_o,\t/a/MEM_aludat [10]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [10],\t/a/EX_regdat2 [10]}),
    .mi({open_n21707,\t/a/EX_regdat2 [10]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [10],_al_u2069_o}),
    .q({\t/a/EX_regdat2 [10],\t/a/MEM_regdat2 [10]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b11|t/a/ex_mem/reg1_b11  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1668_o,\t/a/alu_B_select [1]}),
    .c({_al_u1678_o,\t/a/MEM_aludat [11]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [11],\t/a/EX_regdat2 [11]}),
    .mi({open_n21722,\t/a/EX_regdat2 [11]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [11],_al_u2066_o}),
    .q({\t/a/EX_regdat2 [11],\t/a/MEM_regdat2 [11]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b12|t/a/ex_mem/reg1_b12  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1647_o,\t/a/alu_B_select [1]}),
    .c({_al_u1657_o,\t/a/MEM_aludat [12]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [12],\t/a/EX_regdat2 [12]}),
    .mi({open_n21730,\t/a/EX_regdat2 [12]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [12],_al_u2063_o}),
    .q({\t/a/EX_regdat2 [12],\t/a/MEM_regdat2 [12]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b13|t/a/ex_mem/reg1_b13  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1626_o,\t/a/alu_B_select [1]}),
    .c({_al_u1636_o,\t/a/MEM_aludat [13]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [13],\t/a/EX_regdat2 [13]}),
    .mi({open_n21749,\t/a/EX_regdat2 [13]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [13],_al_u2060_o}),
    .q({\t/a/EX_regdat2 [13],\t/a/MEM_regdat2 [13]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b14|t/a/ex_mem/reg1_b14  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1605_o,\t/a/alu_B_select [1]}),
    .c({_al_u1615_o,\t/a/MEM_aludat [14]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [14],\t/a/EX_regdat2 [14]}),
    .mi({open_n21775,\t/a/EX_regdat2 [14]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [14],_al_u2057_o}),
    .q({\t/a/EX_regdat2 [14],\t/a/MEM_regdat2 [14]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b15|t/a/ex_mem/reg1_b15  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1584_o,\t/a/alu_B_select [1]}),
    .c({_al_u1594_o,\t/a/MEM_aludat [15]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [15],\t/a/EX_regdat2 [15]}),
    .mi({open_n21790,\t/a/EX_regdat2 [15]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [15],_al_u2054_o}),
    .q({\t/a/EX_regdat2 [15],\t/a/MEM_regdat2 [15]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b16|t/a/ex_mem/reg1_b16  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1563_o,\t/a/alu_B_select [1]}),
    .c({_al_u1573_o,\t/a/MEM_aludat [16]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [16],\t/a/EX_regdat2 [16]}),
    .mi({open_n21798,\t/a/EX_regdat2 [16]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [16],_al_u2051_o}),
    .q({\t/a/EX_regdat2 [16],\t/a/MEM_regdat2 [16]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b17|t/a/ex_mem/reg1_b17  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1542_o,\t/a/alu_B_select [1]}),
    .c({_al_u1552_o,\t/a/MEM_aludat [17]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [17],\t/a/EX_regdat2 [17]}),
    .mi({open_n21817,\t/a/EX_regdat2 [17]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [17],_al_u2048_o}),
    .q({\t/a/EX_regdat2 [17],\t/a/MEM_regdat2 [17]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b18|t/a/ex_mem/reg1_b18  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1521_o,\t/a/alu_B_select [1]}),
    .c({_al_u1531_o,\t/a/MEM_aludat [18]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [18],\t/a/EX_regdat2 [18]}),
    .mi({open_n21843,\t/a/EX_regdat2 [18]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [18],_al_u2045_o}),
    .q({\t/a/EX_regdat2 [18],\t/a/MEM_regdat2 [18]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b19|t/a/ex_mem/reg1_b19  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1500_o,\t/a/alu_B_select [1]}),
    .c({_al_u1510_o,\t/a/MEM_aludat [19]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [19],\t/a/EX_regdat2 [19]}),
    .mi({open_n21858,\t/a/EX_regdat2 [19]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [19],_al_u2042_o}),
    .q({\t/a/EX_regdat2 [19],\t/a/MEM_regdat2 [19]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b1|t/a/ex_mem/reg1_b1  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1479_o,\t/a/alu_B_select [1]}),
    .c({_al_u1489_o,\t/a/MEM_aludat [1]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [1],\t/a/EX_regdat2 [1]}),
    .mi({open_n21866,\t/a/EX_regdat2 [1]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [1],_al_u2072_o}),
    .q({\t/a/EX_regdat2 [1],\t/a/MEM_regdat2 [1]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b20|t/a/ex_mem/reg1_b20  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1458_o,\t/a/alu_B_select [1]}),
    .c({_al_u1468_o,\t/a/MEM_aludat [20]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [20],\t/a/EX_regdat2 [20]}),
    .mi({open_n21885,\t/a/EX_regdat2 [20]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [20],_al_u2039_o}),
    .q({\t/a/EX_regdat2 [20],\t/a/MEM_regdat2 [20]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b21|t/a/ex_mem/reg1_b21  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1437_o,\t/a/alu_B_select [1]}),
    .c({_al_u1447_o,\t/a/MEM_aludat [21]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [21],\t/a/EX_regdat2 [21]}),
    .mi({open_n21904,\t/a/EX_regdat2 [21]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [21],_al_u2036_o}),
    .q({\t/a/EX_regdat2 [21],\t/a/MEM_regdat2 [21]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b22|t/a/ex_mem/reg1_b22  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1416_o,\t/a/alu_B_select [1]}),
    .c({_al_u1426_o,\t/a/MEM_aludat [22]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [22],\t/a/EX_regdat2 [22]}),
    .mi({open_n21930,\t/a/EX_regdat2 [22]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [22],_al_u2033_o}),
    .q({\t/a/EX_regdat2 [22],\t/a/MEM_regdat2 [22]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b23|t/a/ex_mem/reg1_b23  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1395_o,\t/a/alu_B_select [1]}),
    .c({_al_u1405_o,\t/a/MEM_aludat [23]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [23],\t/a/EX_regdat2 [23]}),
    .mi({open_n21945,\t/a/EX_regdat2 [23]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [23],_al_u2030_o}),
    .q({\t/a/EX_regdat2 [23],\t/a/MEM_regdat2 [23]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b24|t/a/ex_mem/reg1_b24  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1374_o,\t/a/alu_B_select [1]}),
    .c({_al_u1384_o,\t/a/MEM_aludat [24]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [24],\t/a/EX_regdat2 [24]}),
    .mi({open_n21953,\t/a/EX_regdat2 [24]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [24],_al_u2027_o}),
    .q({\t/a/EX_regdat2 [24],\t/a/MEM_regdat2 [24]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b25|t/a/ex_mem/reg1_b25  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1353_o,\t/a/alu_B_select [1]}),
    .c({_al_u1363_o,\t/a/MEM_aludat [25]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [25],\t/a/EX_regdat2 [25]}),
    .mi({open_n21972,\t/a/EX_regdat2 [25]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [25],_al_u2024_o}),
    .q({\t/a/EX_regdat2 [25],\t/a/MEM_regdat2 [25]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b26|t/a/ex_mem/reg1_b26  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1332_o,\t/a/alu_B_select [1]}),
    .c({_al_u1342_o,\t/a/MEM_aludat [26]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [26],\t/a/EX_regdat2 [26]}),
    .mi({open_n21998,\t/a/EX_regdat2 [26]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [26],_al_u2021_o}),
    .q({\t/a/EX_regdat2 [26],\t/a/MEM_regdat2 [26]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b27|t/a/ex_mem/reg1_b27  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1311_o,\t/a/alu_B_select [1]}),
    .c({_al_u1321_o,\t/a/MEM_aludat [27]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [27],\t/a/EX_regdat2 [27]}),
    .mi({open_n22013,\t/a/EX_regdat2 [27]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [27],_al_u2018_o}),
    .q({\t/a/EX_regdat2 [27],\t/a/MEM_regdat2 [27]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b28|t/a/ex_mem/reg1_b28  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1290_o,\t/a/alu_B_select [1]}),
    .c({_al_u1300_o,\t/a/MEM_aludat [28]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [28],\t/a/EX_regdat2 [28]}),
    .mi({open_n22021,\t/a/EX_regdat2 [28]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [28],_al_u2015_o}),
    .q({\t/a/EX_regdat2 [28],\t/a/MEM_regdat2 [28]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b29|t/a/ex_mem/reg1_b29  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1269_o,\t/a/alu_B_select [1]}),
    .c({_al_u1279_o,\t/a/MEM_aludat [29]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [29],\t/a/EX_regdat2 [29]}),
    .mi({open_n22040,\t/a/EX_regdat2 [29]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [29],_al_u2012_o}),
    .q({\t/a/EX_regdat2 [29],\t/a/MEM_regdat2 [29]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b30|t/a/ex_mem/reg1_b30  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1227_o,\t/a/alu_B_select [1]}),
    .c({_al_u1237_o,\t/a/MEM_aludat [30]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [30],\t/a/EX_regdat2 [30]}),
    .mi({open_n22066,\t/a/EX_regdat2 [30]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [30],_al_u2005_o}),
    .q({\t/a/EX_regdat2 [30],\t/a/MEM_regdat2 [30]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b31|t/a/ex_mem/reg1_b31  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1206_o,\t/a/alu_B_select [1]}),
    .c({_al_u1216_o,\t/a/MEM_aludat [31]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [31],\t/a/EX_regdat2 [31]}),
    .mi({open_n22074,\t/a/EX_regdat2 [31]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [31],_al_u2002_o}),
    .q({\t/a/EX_regdat2 [31],\t/a/MEM_regdat2 [31]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b3|t/a/ex_mem/reg1_b3  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1185_o,\t/a/alu_B_select [1]}),
    .c({_al_u1195_o,\t/a/MEM_aludat [3]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [3],\t/a/EX_regdat2 [3]}),
    .mi({open_n22100,\t/a/EX_regdat2 [3]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [3],_al_u2009_o}),
    .q({\t/a/EX_regdat2 [3],\t/a/MEM_regdat2 [3]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b4|t/a/ex_mem/reg1_b4  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1164_o,\t/a/alu_B_select [1]}),
    .c({_al_u1174_o,\t/a/MEM_aludat [4]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [4],\t/a/EX_regdat2 [4]}),
    .mi({open_n22108,\t/a/EX_regdat2 [4]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [4],_al_u1999_o}),
    .q({\t/a/EX_regdat2 [4],\t/a/MEM_regdat2 [4]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b5|t/a/ex_mem/reg1_b5  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1143_o,\t/a/alu_B_select [1]}),
    .c({_al_u1153_o,\t/a/MEM_aludat [5]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [5],\t/a/EX_regdat2 [5]}),
    .mi({open_n22134,\t/a/EX_regdat2 [5]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [5],_al_u1996_o}),
    .q({\t/a/EX_regdat2 [5],\t/a/MEM_regdat2 [5]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b6|t/a/ex_mem/reg1_b6  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1122_o,\t/a/alu_B_select [1]}),
    .c({_al_u1132_o,\t/a/MEM_aludat [6]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [6],\t/a/EX_regdat2 [6]}),
    .mi({open_n22149,\t/a/EX_regdat2 [6]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [6],_al_u1993_o}),
    .q({\t/a/EX_regdat2 [6],\t/a/MEM_regdat2 [6]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b7|t/a/ex_mem/reg1_b7  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1101_o,\t/a/alu_B_select [1]}),
    .c({_al_u1111_o,\t/a/MEM_aludat [7]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [7],\t/a/EX_regdat2 [7]}),
    .mi({open_n22157,\t/a/EX_regdat2 [7]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [7],_al_u1990_o}),
    .q({\t/a/EX_regdat2 [7],\t/a/MEM_regdat2 [7]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTF1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUTG0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUTG1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000010011),
    .INIT_LUTF1(16'b1010101100000001),
    .INIT_LUTG0(16'b0000001000010011),
    .INIT_LUTG1(16'b1010101100000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b8|t/a/ex_mem/reg1_b8  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1080_o,\t/a/alu_B_select [1]}),
    .c({_al_u1090_o,\t/a/MEM_aludat [8]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [8],\t/a/EX_regdat2 [8]}),
    .mi({open_n22176,\t/a/EX_regdat2 [8]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [8],_al_u1987_o}),
    .q({\t/a/EX_regdat2 [8],\t/a/MEM_regdat2 [8]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg0_b9|t/a/ex_mem/reg1_b9  (
    .a({_al_u1049_o,\t/a/alu_B_select [0]}),
    .b({_al_u1059_o,\t/a/alu_B_select [1]}),
    .c({_al_u1069_o,\t/a/MEM_aludat [9]}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [9],\t/a/EX_regdat2 [9]}),
    .mi({open_n22202,\t/a/EX_regdat2 [9]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat2 [9],_al_u1979_o}),
    .q({\t/a/EX_regdat2 [9],\t/a/MEM_regdat2 [9]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(0*(C@(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTF1("(~0*~D*(C@(B*A)))"),
    //.LUTG0("(1*(C@(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D)))"),
    //.LUTG1("(~1*~D*(C@(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000001111000),
    .INIT_LUTG0(16'b0011110001011010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg1_b0|t/a/id_ex/reg1_b1  (
    .a({_al_u2777_o,\t/a/condition/n9 }),
    .b({_al_u2790_o,\t/a/condition/n10 }),
    .c({\t/a/ID_fun3 [0],\t/a/ID_fun3 [0]}),
    .clk(clock_pad),
    .d({\t/a/ID_fun3 [1],\t/a/ID_fun3 [1]}),
    .e({\t/a/ID_fun3 [2],\t/a/ID_fun3 [2]}),
    .mi({\t/a/ID_fun3 [0],\t/a/ID_fun3 [1]}),
    .sr(rst_pad),
    .f({_al_u2791_o,_al_u2766_o}),
    .q({\t/a/EX_fun3 [0],\t/a/EX_fun3 [1]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(D*C)*~(0*A))"),
    //.LUTF1("~(~B*~A*~(D*C))"),
    //.LUTG0("(~B*~(D*C)*~(1*A))"),
    //.LUTG1("~(~B*~A*~(D*C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100110011),
    .INIT_LUTF1(16'b1111111011101110),
    .INIT_LUTG0(16'b0000000100010001),
    .INIT_LUTG1(16'b1111111011101110),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg3_b2|t/a/ex_mem/reg0_b2  (
    .a({\t/a/aluin/sel1_b22/B9 ,\t/a/aluin/n12_lutinv }),
    .b({_al_u2007_o,_al_u1802_o}),
    .c({_al_u1803_o,_al_u1984_o}),
    .clk(clock_pad),
    .d({\t/a/EX_rs2 [2],\t/a/EX_rs2 [2]}),
    .e({open_n22223,\t/a/EX_rd [2]}),
    .mi({\t/a/ID_rs2 [2],\t/a/EX_rd [2]}),
    .sr(rst_pad),
    .f({\t/a/EX_B [22],_al_u2093_o}),
    .q({\t/a/EX_rs2 [2],\t/a/MEM_rd [2]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(71)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("((C@B)*(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0001010000101000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg5_b0|t/a/if_id/reg2_b0  (
    .a({_al_u2111_o,\t/a/if_id/n9 }),
    .b({_al_u2119_o,\t/busarbitration/n3 }),
    .c({\t/a/ID_rd [0],\t/busarbitration/instruction [7]}),
    .clk(clock_pad),
    .d({\t/a/ID_rd [4],i_data[7]}),
    .mi({\t/a/ID_rd [0],open_n22250}),
    .sr(rst_pad),
    .f({_al_u2806_o,open_n22251}),
    .q({\t/a/EX_rd [0],\t/a/ID_rd [0]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg5_b3|t/a/if_id/reg2_b3  (
    .a({open_n22255,\t/a/if_id/n9 }),
    .b({open_n22256,\t/busarbitration/n3 }),
    .c({\t/a/ID_rd [3],\t/busarbitration/instruction [10]}),
    .clk(clock_pad),
    .d({_al_u2113_o,i_data[10]}),
    .mi({\t/a/ID_rd [3],open_n22268}),
    .sr(rst_pad),
    .f({_al_u2799_o,open_n22269}),
    .q({\t/a/EX_rd [3],\t/a/ID_rd [3]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("((C@B)*(D@A))"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("((C@B)*(D@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0001010000101000),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0001010000101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg5_b4|t/a/if_id/reg2_b4  (
    .a({_al_u1956_o,\t/a/if_id/n9 }),
    .b({_al_u1960_o,\t/busarbitration/n3 }),
    .c({\t/a/ID_rd [2],\t/busarbitration/instruction [11]}),
    .clk(clock_pad),
    .d({\t/a/ID_rd [4],i_data[11]}),
    .mi({\t/a/ID_rd [4],open_n22277}),
    .sr(rst_pad),
    .f({_al_u2793_o,open_n22289}),
    .q({\t/a/EX_rd [4],\t/a/ID_rd [4]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0101010000010000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0101010000010000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg6_b0|t/a/if_id/reg6_b0  (
    .a({_al_u2803_o,\t/a/if_id/n9 }),
    .b({\t/a/ID_op [0],\t/busarbitration/n3 }),
    .c({\t/a/ID_op [1],\t/busarbitration/instruction [0]}),
    .clk(clock_pad),
    .d({\t/a/ID_op [2],i_data[0]}),
    .mi({\t/a/ID_op [0],open_n22297}),
    .sr(rst_pad),
    .f({\t/a/n0_lutinv ,open_n22309}),
    .q({\t/a/EX_op [0],\t/a/ID_op [0]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg6_b2|t/a/if_id/reg6_b2  (
    .a({_al_u1747_o,open_n22313}),
    .b({\t/a/ID_op [0],open_n22314}),
    .c({\t/a/ID_op [1],\t/instruction$2$_neg_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_op [2],\t/a/if_id/n9 }),
    .mi({\t/a/ID_op [2],open_n22319}),
    .sr(rst_pad),
    .f({\t/a/condition/n1_lutinv ,open_n22331}),
    .q({\t/a/EX_op [2],\t/a/ID_op [2]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg6_b3|t/a/if_id/reg6_b6  (
    .a({\t/a/ID_op [3],\t/a/if_id/n9 }),
    .b({\t/a/ID_op [4],\t/busarbitration/n3 }),
    .c({\t/a/ID_op [5],\t/busarbitration/instruction [6]}),
    .clk(clock_pad),
    .d({\t/a/ID_op [6],i_data[6]}),
    .mi({\t/a/ID_op [3],open_n22346}),
    .sr(rst_pad),
    .f({_al_u2803_o,open_n22347}),
    .q({\t/a/EX_op [3],\t/a/ID_op [6]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(D*C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101010000010000),
    .INIT_LUT1(16'b0001000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg6_b4|t/a/if_id/reg6_b5  (
    .a({\t/a/ID_op [3],\t/a/if_id/n9 }),
    .b({\t/a/ID_op [4],\t/busarbitration/n3 }),
    .c({\t/a/ID_op [5],\t/busarbitration/instruction [5]}),
    .clk(clock_pad),
    .d({\t/a/ID_op [6],i_data[5]}),
    .mi({\t/a/ID_op [4],open_n22362}),
    .sr(rst_pad),
    .f({_al_u1747_o,open_n22363}),
    .q({\t/a/EX_op [4],\t/a/ID_op [5]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0*D))"),
    //.LUTF1("(C*B*A*~(0*D))"),
    //.LUTG0("(C*B*A*~(1*D))"),
    //.LUTG1("(C*B*A*~(1*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000010000000),
    .INIT_LUTF1(16'b1000000010000000),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg6_b5|t/a/ex_mem/reg2_b5  (
    .a({_al_u2608_o,_al_u2608_o}),
    .b({\t/a/risk_jump/n35_lutinv ,\t/a/risk_jump/n11_lutinv }),
    .c({\t/a/condition/n1_lutinv ,\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({_al_u1740_o,_al_u1740_o}),
    .e({\t/a/EX_op [5],\t/a/EX_op [5]}),
    .mi({\t/a/ID_op [5],\t/a/EX_op [5]}),
    .sr(rst_pad),
    .f({_al_u2609_o,_al_u2615_o}),
    .q({\t/a/EX_op [5],\t/a/MEM_op [5]}));  // flow_line_reg.v(191)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUT1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111100010),
    .INIT_LUT1(16'b1111001111100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b11|t/a/id_ex/reg7_b30  (
    .a({_al_u2807_o,_al_u2807_o}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/ID_memstraddr [11],\t/a/ID_memstraddr [30]}),
    .clk(clock_pad),
    .d({\t/memstraddress [11],\t/memstraddress [30]}),
    .mi({\t/a/ID_memstraddr [11],\t/a/ID_memstraddr [30]}),
    .sr(rst_pad),
    .f({_al_u2883_o,_al_u2829_o}),
    .q({\t/a/EX_memstraddr [11],\t/a/EX_memstraddr [30]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTF1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTG0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTG1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111100010),
    .INIT_LUTF1(16'b1111001111100010),
    .INIT_LUTG0(16'b1111001111100010),
    .INIT_LUTG1(16'b1111001111100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b13|t/a/id_ex/reg7_b29  (
    .a({_al_u2807_o,_al_u2807_o}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/ID_memstraddr [13],\t/a/ID_memstraddr [29]}),
    .clk(clock_pad),
    .d({\t/memstraddress [13],\t/memstraddress [29]}),
    .mi({\t/a/ID_memstraddr [13],\t/a/ID_memstraddr [29]}),
    .sr(rst_pad),
    .f({_al_u2878_o,_al_u2834_o}),
    .q({\t/a/EX_memstraddr [13],\t/a/EX_memstraddr [29]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTF1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTG0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTG1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111100010),
    .INIT_LUTF1(16'b1111001111100010),
    .INIT_LUTG0(16'b1111001111100010),
    .INIT_LUTG1(16'b1111001111100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b14|t/a/id_ex/reg7_b26  (
    .a({_al_u2807_o,_al_u2807_o}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/ID_memstraddr [14],\t/a/ID_memstraddr [26]}),
    .clk(clock_pad),
    .d({\t/memstraddress [14],\t/memstraddress [26]}),
    .mi({\t/a/ID_memstraddr [14],\t/a/ID_memstraddr [26]}),
    .sr(rst_pad),
    .f({_al_u2875_o,_al_u2841_o}),
    .q({\t/a/EX_memstraddr [14],\t/a/EX_memstraddr [26]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUT1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111100010),
    .INIT_LUT1(16'b1111001111100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b15|t/a/id_ex/reg7_b25  (
    .a({_al_u2807_o,_al_u2807_o}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/ID_memstraddr [15],\t/a/ID_memstraddr [25]}),
    .clk(clock_pad),
    .d({\t/memstraddress [15],\t/memstraddress [25]}),
    .mi({\t/a/ID_memstraddr [15],\t/a/ID_memstraddr [25]}),
    .sr(rst_pad),
    .f({_al_u2872_o,_al_u2844_o}),
    .q({\t/a/EX_memstraddr [15],\t/a/EX_memstraddr [25]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUT1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111001111100010),
    .INIT_LUT1(16'b1111001111100010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b16|t/a/id_ex/reg7_b24  (
    .a({_al_u2807_o,_al_u2807_o}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/ID_memstraddr [16],\t/a/ID_memstraddr [24]}),
    .clk(clock_pad),
    .d({\t/memstraddress [16],\t/memstraddress [24]}),
    .mi({\t/a/ID_memstraddr [16],\t/a/ID_memstraddr [24]}),
    .sr(rst_pad),
    .f({_al_u2869_o,_al_u2847_o}),
    .q({\t/a/EX_memstraddr [16],\t/a/EX_memstraddr [24]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTF1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTG0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTG1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111100010),
    .INIT_LUTF1(16'b1111001111100010),
    .INIT_LUTG0(16'b1111001111100010),
    .INIT_LUTG1(16'b1111001111100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b1|t/a/id_ex/reg7_b23  (
    .a({_al_u2807_o,_al_u2807_o}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/ID_memstraddr [1],\t/a/ID_memstraddr [23]}),
    .clk(clock_pad),
    .d({\t/memstraddress [1],\t/memstraddress [23]}),
    .mi({\t/a/ID_memstraddr [1],\t/a/ID_memstraddr [23]}),
    .sr(rst_pad),
    .f({_al_u2888_o,_al_u2850_o}),
    .q({\t/a/EX_memstraddr [1],\t/a/EX_memstraddr [23]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_LSLICE #(
    //.LUTF0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTF1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTG0("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    //.LUTG1("(~(~D*~A)*~(C)*~(B)+~(~D*~A)*C*~(B)+~(~(~D*~A))*C*B+~(~D*~A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001111100010),
    .INIT_LUTF1(16'b1111001111100010),
    .INIT_LUTG0(16'b1111001111100010),
    .INIT_LUTG1(16'b1111001111100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg7_b2|t/a/id_ex/reg7_b20  (
    .a({_al_u2807_o,_al_u2807_o}),
    .b({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .c({\t/a/ID_memstraddr [2],\t/a/ID_memstraddr [20]}),
    .clk(clock_pad),
    .d({\t/memstraddress [2],\t/memstraddress [20]}),
    .mi({\t/a/ID_memstraddr [2],\t/a/ID_memstraddr [20]}),
    .sr(rst_pad),
    .f({_al_u2860_o,_al_u2857_o}),
    .q({\t/a/EX_memstraddr [2],\t/a/EX_memstraddr [20]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b0|t/a/id_ex/reg8_b9  (
    .a({_al_u333_o,_al_u333_o}),
    .b({_al_u994_o,_al_u343_o}),
    .c({_al_u1004_o,_al_u353_o}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [0],\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [0],\t/a/ID_read_dat1 [9]}),
    .q({\t/a/EX_regdat1 [0],\t/a/EX_regdat1 [9]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b10|t/a/id_ex/reg8_b30  (
    .a({_al_u333_o,_al_u333_o}),
    .b({_al_u973_o,_al_u511_o}),
    .c({_al_u983_o,_al_u521_o}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [10],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [10],\t/a/ID_read_dat1 [30]}),
    .q({\t/a/EX_regdat1 [10],\t/a/EX_regdat1 [30]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b11|t/a/id_ex/reg8_b27  (
    .a({_al_u333_o,_al_u333_o}),
    .b({_al_u952_o,_al_u595_o}),
    .c({_al_u962_o,_al_u605_o}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [11],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [11],\t/a/ID_read_dat1 [27]}),
    .q({\t/a/EX_regdat1 [11],\t/a/EX_regdat1 [27]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b12|t/a/id_ex/reg8_b26  (
    .a({_al_u333_o,_al_u333_o}),
    .b({_al_u931_o,_al_u616_o}),
    .c({_al_u941_o,_al_u626_o}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [12],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [12],\t/a/ID_read_dat1 [26]}),
    .q({\t/a/EX_regdat1 [12],\t/a/EX_regdat1 [26]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b13|t/a/id_ex/reg8_b23  (
    .a({_al_u333_o,_al_u333_o}),
    .b({_al_u910_o,_al_u679_o}),
    .c({_al_u920_o,_al_u689_o}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [13],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [13],\t/a/ID_read_dat1 [23]}),
    .q({\t/a/EX_regdat1 [13],\t/a/EX_regdat1 [23]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b14|t/a/id_ex/reg8_b22  (
    .a({_al_u333_o,_al_u333_o}),
    .b({_al_u889_o,_al_u700_o}),
    .c({_al_u899_o,_al_u710_o}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [14],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [14],\t/a/ID_read_dat1 [22]}),
    .q({\t/a/EX_regdat1 [14],\t/a/EX_regdat1 [22]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  EG_PHY_MSLICE #(
    //.LUT0("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    //.LUT1("((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010101100000001),
    .INIT_LUT1(16'b1010101100000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/id_ex/reg8_b15|t/a/id_ex/reg8_b19  (
    .a({_al_u333_o,_al_u333_o}),
    .b({_al_u868_o,_al_u784_o}),
    .c({_al_u878_o,_al_u794_o}),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [15],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({\t/a/ID_read_dat1 [15],\t/a/ID_read_dat1 [19]}),
    .q({\t/a/EX_regdat1 [15],\t/a/EX_regdat1 [19]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0101010000010000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0101010000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b0|t/a/id_ex/reg2_b0  (
    .a({\t/a/if_id/n9 ,\t/a/condition/n5 [5]}),
    .b({\t/busarbitration/n3 ,\t/a/condition/n0_lutinv }),
    .c({\t/busarbitration/instruction [25],\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({i_data[25],\t/a/condition/sel1/B2 }),
    .e({open_n22610,\t/a/ID_fun7 [0]}),
    .mi({open_n22612,\t/a/ID_fun7 [0]}),
    .sr(rst_pad),
    .f({open_n22624,\t/a/ID_jump_addr [5]}),
    .q({\t/a/ID_fun7 [0],\t/a/EX_fun7 [0]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0101010000010000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0101010000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b1|t/a/id_ex/reg2_b1  (
    .a({\t/a/if_id/n9 ,\t/a/condition/n5 [6]}),
    .b({\t/busarbitration/n3 ,\t/a/condition/n0_lutinv }),
    .c({\t/busarbitration/instruction [26],\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({i_data[26],\t/a/condition/sel1/B2 }),
    .e({open_n22629,\t/a/ID_fun7 [1]}),
    .mi({open_n22631,\t/a/ID_fun7 [1]}),
    .sr(rst_pad),
    .f({open_n22643,\t/a/ID_jump_addr [6]}),
    .q({\t/a/ID_fun7 [1],\t/a/EX_fun7 [1]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0101010000010000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0101010000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b2|t/a/id_ex/reg2_b2  (
    .a({\t/a/if_id/n9 ,\t/a/condition/n5 [7]}),
    .b({\t/busarbitration/n3 ,\t/a/condition/n0_lutinv }),
    .c({\t/busarbitration/instruction [27],\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({i_data[27],\t/a/condition/sel1/B2 }),
    .e({open_n22648,\t/a/ID_fun7 [2]}),
    .mi({open_n22650,\t/a/ID_fun7 [2]}),
    .sr(rst_pad),
    .f({open_n22662,\t/a/ID_jump_addr [7]}),
    .q({\t/a/ID_fun7 [2],\t/a/EX_fun7 [2]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0101010000010000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0101010000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b3|t/a/id_ex/reg2_b3  (
    .a({\t/a/if_id/n9 ,\t/a/condition/n5 [8]}),
    .b({\t/busarbitration/n3 ,\t/a/condition/n0_lutinv }),
    .c({\t/busarbitration/instruction [28],\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({i_data[28],\t/a/condition/sel1/B2 }),
    .e({open_n22667,\t/a/ID_fun7 [3]}),
    .mi({open_n22669,\t/a/ID_fun7 [3]}),
    .sr(rst_pad),
    .f({open_n22681,\t/a/ID_jump_addr [8]}),
    .q({\t/a/ID_fun7 [3],\t/a/EX_fun7 [3]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0101010000010000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0101010000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b4|t/a/id_ex/reg2_b4  (
    .a({\t/a/if_id/n9 ,\t/a/condition/n5 [9]}),
    .b({\t/busarbitration/n3 ,\t/a/condition/n0_lutinv }),
    .c({\t/busarbitration/instruction [29],\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({i_data[29],\t/a/condition/sel1/B2 }),
    .e({open_n22686,\t/a/ID_fun7 [4]}),
    .mi({open_n22688,\t/a/ID_fun7 [4]}),
    .sr(rst_pad),
    .f({open_n22700,\t/a/ID_jump_addr [9]}),
    .q({\t/a/ID_fun7 [4],\t/a/EX_fun7 [4]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(139)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(~B*~(~(0*C)*~(D*A)))"),
    //.LUTF1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~B*~(~(1*C)*~(D*A)))"),
    //.LUTG1("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001000000000),
    .INIT_LUTF1(16'b0101010000010000),
    .INIT_LUTG0(16'b0011001000110000),
    .INIT_LUTG1(16'b0101010000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg1_b5|t/a/id_ex/reg2_b5  (
    .a({\t/a/if_id/n9 ,\t/a/condition/n5 [10]}),
    .b({\t/busarbitration/n3 ,\t/a/condition/n0_lutinv }),
    .c({\t/busarbitration/instruction [30],\t/a/condition/n1_lutinv }),
    .clk(clock_pad),
    .d({i_data[30],\t/a/condition/sel1/B2 }),
    .e({open_n22705,\t/a/ID_fun7 [5]}),
    .mi({open_n22707,\t/a/ID_fun7 [5]}),
    .sr(rst_pad),
    .f({open_n22719,\t/a/ID_jump_addr [10]}),
    .q({\t/a/ID_fun7 [5],\t/a/EX_fun7 [5]}));  // flow_line_reg.v(139)
  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b10|t/a/if_id/reg5_b8  (
    .b({\t/a/MEM_aludat [10],\t/a/MEM_aludat [8]}),
    .c({\t/memstraddress [10],\t/memstraddress [8]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .mi({\t/memstraddress [10],\t/memstraddress [8]}),
    .sr(rst_pad),
    .f({addr[10],addr[8]}),
    .q({\t/a/ID_memstraddr [10],\t/a/ID_memstraddr [8]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b11|t/a/if_id/reg5_b30  (
    .b({\t/a/MEM_aludat [11],\t/a/MEM_aludat [30]}),
    .c({\t/memstraddress [11],\t/memstraddress [30]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .mi({\t/memstraddress [11],\t/memstraddress [30]}),
    .sr(rst_pad),
    .f({addr[11],addr[30]}),
    .q({\t/a/ID_memstraddr [11],\t/a/ID_memstraddr [30]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b12|t/a/if_id/reg5_b28  (
    .b({\t/a/MEM_aludat [12],\t/a/MEM_aludat [28]}),
    .c({\t/memstraddress [12],\t/memstraddress [28]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .mi({\t/memstraddress [12],\t/memstraddress [28]}),
    .sr(rst_pad),
    .f({addr[12],addr[28]}),
    .q({\t/a/ID_memstraddr [12],\t/a/ID_memstraddr [28]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b13|t/a/if_id/reg5_b27  (
    .b({\t/a/MEM_aludat [13],\t/a/MEM_aludat [27]}),
    .c({\t/memstraddress [13],\t/memstraddress [27]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .mi({\t/memstraddress [13],\t/memstraddress [27]}),
    .sr(rst_pad),
    .f({addr[13],addr[27]}),
    .q({\t/a/ID_memstraddr [13],\t/a/ID_memstraddr [27]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b14|t/a/if_id/reg5_b25  (
    .b({\t/a/MEM_aludat [14],\t/a/MEM_aludat [25]}),
    .c({\t/memstraddress [14],\t/memstraddress [25]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .mi({\t/memstraddress [14],\t/memstraddress [25]}),
    .sr(rst_pad),
    .f({addr[14],addr[25]}),
    .q({\t/a/ID_memstraddr [14],\t/a/ID_memstraddr [25]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b15|t/a/if_id/reg5_b23  (
    .b({\t/a/MEM_aludat [15],\t/a/MEM_aludat [23]}),
    .c({\t/memstraddress [15],\t/memstraddress [23]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .mi({\t/memstraddress [15],\t/memstraddress [23]}),
    .sr(rst_pad),
    .f({addr[15],addr[23]}),
    .q({\t/a/ID_memstraddr [15],\t/a/ID_memstraddr [23]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b16|t/a/if_id/reg5_b21  (
    .b({\t/a/MEM_aludat [16],\t/a/MEM_aludat [21]}),
    .c({\t/memstraddress [16],\t/memstraddress [21]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .mi({\t/memstraddress [16],\t/memstraddress [21]}),
    .sr(rst_pad),
    .f({addr[16],addr[21]}),
    .q({\t/a/ID_memstraddr [16],\t/a/ID_memstraddr [21]}));  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  // flow_line_reg.v(71)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/if_id/reg5_b17|t/a/if_id/reg5_b20  (
    .b({\t/a/MEM_aludat [17],\t/a/MEM_aludat [20]}),
    .c({\t/memstraddress [17],\t/memstraddress [20]}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/busarbitration/n3 ,\t/busarbitration/n3 }),
    .mi({\t/memstraddress [17],\t/memstraddress [20]}),
    .sr(rst_pad),
    .f({addr[17],addr[20]}),
    .q({\t/a/ID_memstraddr [17],\t/a/ID_memstraddr [20]}));  // flow_line_reg.v(71)
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u11_al_u2955  (
    .a({\t/memstraddress [13],\t/memstraddress [11]}),
    .b({\t/memstraddress [14],\t/memstraddress [12]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [13],\t/a/IF_skip_addr [11]}),
    .e({\t/a/IF_skip_addr [14],\t/a/IF_skip_addr [12]}),
    .fci(\t/a/instr/add0/c11 ),
    .f({\t/a/instr/n12 [13],\t/a/instr/n12 [11]}),
    .fco(\t/a/instr/add0/c15 ),
    .fx({\t/a/instr/n12 [14],\t/a/instr/n12 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u15_al_u2956  (
    .a({\t/memstraddress [17],\t/memstraddress [15]}),
    .b({\t/memstraddress [18],\t/memstraddress [16]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [17],\t/a/IF_skip_addr [15]}),
    .e({\t/a/IF_skip_addr [18],\t/a/IF_skip_addr [16]}),
    .fci(\t/a/instr/add0/c15 ),
    .f({\t/a/instr/n12 [17],\t/a/instr/n12 [15]}),
    .fco(\t/a/instr/add0/c19 ),
    .fx({\t/a/instr/n12 [18],\t/a/instr/n12 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u19_al_u2957  (
    .a({\t/memstraddress [21],\t/memstraddress [19]}),
    .b({\t/memstraddress [22],\t/memstraddress [20]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [21],\t/a/IF_skip_addr [19]}),
    .e({\t/a/IF_skip_addr [22],\t/a/IF_skip_addr [20]}),
    .fci(\t/a/instr/add0/c19 ),
    .f({\t/a/instr/n12 [21],\t/a/instr/n12 [19]}),
    .fco(\t/a/instr/add0/c23 ),
    .fx({\t/a/instr/n12 [22],\t/a/instr/n12 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u23_al_u2958  (
    .a({\t/memstraddress [25],\t/memstraddress [23]}),
    .b({\t/memstraddress [26],\t/memstraddress [24]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [25],\t/a/IF_skip_addr [23]}),
    .e({\t/a/IF_skip_addr [26],\t/a/IF_skip_addr [24]}),
    .fci(\t/a/instr/add0/c23 ),
    .f({\t/a/instr/n12 [25],\t/a/instr/n12 [23]}),
    .fco(\t/a/instr/add0/c27 ),
    .fx({\t/a/instr/n12 [26],\t/a/instr/n12 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u27_al_u2959  (
    .a({\t/memstraddress [29],\t/memstraddress [27]}),
    .b({\t/memstraddress [30],\t/memstraddress [28]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [29],\t/a/IF_skip_addr [27]}),
    .e({\t/a/IF_skip_addr [30],\t/a/IF_skip_addr [28]}),
    .fci(\t/a/instr/add0/c27 ),
    .f({\t/a/instr/n12 [29],\t/a/instr/n12 [27]}),
    .fco(\t/a/instr/add0/c31 ),
    .fx({\t/a/instr/n12 [30],\t/a/instr/n12 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u31_al_u2960  (
    .a({open_n22949,\t/memstraddress [31]}),
    .c(2'b00),
    .d({open_n22954,\t/a/IF_skip_addr [31]}),
    .fci(\t/a/instr/add0/c31 ),
    .f({open_n22971,\t/a/instr/n12 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u3_al_u2953  (
    .a({\t/memstraddress [5],\t/memstraddress [3]}),
    .b({\t/memstraddress [6],\t/memstraddress [4]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [5],\t/a/IF_skip_addr [3]}),
    .e({\t/a/IF_skip_addr [6],\t/a/IF_skip_addr [4]}),
    .fci(\t/a/instr/add0/c3 ),
    .f({\t/a/instr/n12 [5],\t/a/instr/n12 [3]}),
    .fco(\t/a/instr/add0/c7 ),
    .fx({\t/a/instr/n12 [6],\t/a/instr/n12 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add0/u7_al_u2954  (
    .a({\t/memstraddress [9],\t/memstraddress [7]}),
    .b({\t/memstraddress [10],\t/memstraddress [8]}),
    .c(2'b00),
    .d({\t/a/IF_skip_addr [9],\t/a/IF_skip_addr [7]}),
    .e({\t/a/IF_skip_addr [10],\t/a/IF_skip_addr [8]}),
    .fci(\t/a/instr/add0/c7 ),
    .f({\t/a/instr/n12 [9],\t/a/instr/n12 [7]}),
    .fco(\t/a/instr/add0/c11 ),
    .fx({\t/a/instr/n12 [10],\t/a/instr/n12 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add0/ucin_al_u2952"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/add0/ucin_al_u2952  (
    .a({\t/memstraddress [1],1'b0}),
    .b({\t/memstraddress [2],\t/memstraddress [0]}),
    .c(2'b00),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({\t/a/IF_skip_addr [1],1'b1}),
    .e({\t/a/IF_skip_addr [2],1'b0}),
    .mi({open_n23014,\t/memstraddress [0]}),
    .sr(rst_pad),
    .f({\t/a/instr/n12 [1],open_n23026}),
    .fco(\t/a/instr/add0/c3 ),
    .fx({\t/a/instr/n12 [2],\t/a/instr/n12 [0]}),
    .q({open_n23027,\t/a/ID_memstraddr [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u11_al_u2972  (
    .a({\t/memstraddress [15],\t/memstraddress [13]}),
    .b({\t/memstraddress [16],\t/memstraddress [14]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c11 ),
    .f({\t/a/instr/n16 [13],\t/a/instr/n16 [11]}),
    .fco(\t/a/instr/add2/c15 ),
    .fx({\t/a/instr/n16 [14],\t/a/instr/n16 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u15_al_u2973  (
    .a({\t/memstraddress [19],\t/memstraddress [17]}),
    .b({\t/memstraddress [20],\t/memstraddress [18]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c15 ),
    .f({\t/a/instr/n16 [17],\t/a/instr/n16 [15]}),
    .fco(\t/a/instr/add2/c19 ),
    .fx({\t/a/instr/n16 [18],\t/a/instr/n16 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u19_al_u2974  (
    .a({\t/memstraddress [23],\t/memstraddress [21]}),
    .b({\t/memstraddress [24],\t/memstraddress [22]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c19 ),
    .f({\t/a/instr/n16 [21],\t/a/instr/n16 [19]}),
    .fco(\t/a/instr/add2/c23 ),
    .fx({\t/a/instr/n16 [22],\t/a/instr/n16 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u23_al_u2975  (
    .a({\t/memstraddress [27],\t/memstraddress [25]}),
    .b({\t/memstraddress [28],\t/memstraddress [26]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c23 ),
    .f({\t/a/instr/n16 [25],\t/a/instr/n16 [23]}),
    .fco(\t/a/instr/add2/c27 ),
    .fx({\t/a/instr/n16 [26],\t/a/instr/n16 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u27_al_u2976  (
    .a({\t/memstraddress [31],\t/memstraddress [29]}),
    .b({open_n23100,\t/memstraddress [30]}),
    .c(2'b00),
    .d(2'b00),
    .e({open_n23103,1'b0}),
    .fci(\t/a/instr/add2/c27 ),
    .f({\t/a/instr/n16 [29],\t/a/instr/n16 [27]}),
    .fx({open_n23119,\t/a/instr/n16 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u3_al_u2970  (
    .a({\t/memstraddress [7],\t/memstraddress [5]}),
    .b({\t/memstraddress [8],\t/memstraddress [6]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c3 ),
    .f({\t/a/instr/n16 [5],\t/a/instr/n16 [3]}),
    .fco(\t/a/instr/add2/c7 ),
    .fx({\t/a/instr/n16 [6],\t/a/instr/n16 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \t/a/instr/add2/u7_al_u2971  (
    .a({\t/memstraddress [11],\t/memstraddress [9]}),
    .b({\t/memstraddress [12],\t/memstraddress [10]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\t/a/instr/add2/c7 ),
    .f({\t/a/instr/n16 [9],\t/a/instr/n16 [7]}),
    .fco(\t/a/instr/add2/c11 ),
    .fx({\t/a/instr/n16 [10],\t/a/instr/n16 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("t/a/instr/add2/ucin_al_u2969"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/add2/ucin_al_u2969  (
    .a({\t/memstraddress [3],1'b0}),
    .b({\t/memstraddress [4],\t/memstraddress [2]}),
    .c(2'b00),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d(2'b01),
    .e(2'b01),
    .mi(\t/memstraddress [4:3]),
    .sr(rst_pad),
    .f({\t/a/instr/n16 [1],open_n23170}),
    .fco(\t/a/instr/add2/c3 ),
    .fx({\t/a/instr/n16 [2],\t/a/instr/n16 [0]}),
    .q(\t/a/ID_memstraddr [4:3]));
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b0  (
    .a({_al_u2890_o,_al_u2890_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [0],\t/a/ID_memstraddr [0]}),
    .mi({open_n23182,\t/memstraddress [0]}),
    .sr(rst_pad),
    .q({open_n23188,\t/memstraddress [0]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b1  (
    .a({_al_u2887_o,_al_u2887_o}),
    .b({\t/a/instr/n12 [1],\t/a/instr/n12 [1]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2888_o,_al_u2888_o}),
    .mi({open_n23200,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23206,\t/memstraddress [1]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b10  (
    .a({_al_u2885_o,_al_u2885_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [10],\t/a/ID_memstraddr [10]}),
    .mi({open_n23218,\t/memstraddress [10]}),
    .sr(rst_pad),
    .q({open_n23224,\t/memstraddress [10]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b11  (
    .a({_al_u2882_o,_al_u2882_o}),
    .b({\t/a/instr/n12 [11],\t/a/instr/n12 [11]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2883_o,_al_u2883_o}),
    .mi({open_n23236,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23242,\t/memstraddress [11]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b12  (
    .a({_al_u2880_o,_al_u2880_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [12],\t/a/ID_memstraddr [12]}),
    .mi({open_n23254,\t/memstraddress [12]}),
    .sr(rst_pad),
    .q({open_n23260,\t/memstraddress [12]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b13  (
    .a({_al_u2877_o,_al_u2877_o}),
    .b({\t/a/instr/n12 [13],\t/a/instr/n12 [13]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2878_o,_al_u2878_o}),
    .mi({open_n23272,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23278,\t/memstraddress [13]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b14  (
    .a({_al_u2874_o,_al_u2874_o}),
    .b({\t/a/instr/n12 [14],\t/a/instr/n12 [14]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2875_o,_al_u2875_o}),
    .mi({open_n23290,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23296,\t/memstraddress [14]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b15  (
    .a({_al_u2871_o,_al_u2871_o}),
    .b({\t/a/instr/n12 [15],\t/a/instr/n12 [15]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2872_o,_al_u2872_o}),
    .mi({open_n23308,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23314,\t/memstraddress [15]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b16  (
    .a({_al_u2868_o,_al_u2868_o}),
    .b({\t/a/instr/n12 [16],\t/a/instr/n12 [16]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2869_o,_al_u2869_o}),
    .mi({open_n23326,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23332,\t/memstraddress [16]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b17  (
    .a({_al_u2866_o,_al_u2866_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [17],\t/a/ID_memstraddr [17]}),
    .mi({open_n23344,\t/memstraddress [17]}),
    .sr(rst_pad),
    .q({open_n23350,\t/memstraddress [17]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b18  (
    .a({_al_u2864_o,_al_u2864_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [18],\t/a/ID_memstraddr [18]}),
    .mi({open_n23362,\t/memstraddress [18]}),
    .sr(rst_pad),
    .q({open_n23368,\t/memstraddress [18]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b19  (
    .a({_al_u2862_o,_al_u2862_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [19],\t/a/ID_memstraddr [19]}),
    .mi({open_n23380,\t/memstraddress [19]}),
    .sr(rst_pad),
    .q({open_n23386,\t/memstraddress [19]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("SET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b2  (
    .a({_al_u2859_o,_al_u2859_o}),
    .b({\t/a/instr/n12 [2],\t/a/instr/n12 [2]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2860_o,_al_u2860_o}),
    .mi({open_n23398,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23404,\t/memstraddress [2]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b20  (
    .a({_al_u2856_o,_al_u2856_o}),
    .b({\t/a/instr/n12 [20],\t/a/instr/n12 [20]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2857_o,_al_u2857_o}),
    .mi({open_n23416,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23422,\t/memstraddress [20]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b21  (
    .a({_al_u2854_o,_al_u2854_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [21],\t/a/ID_memstraddr [21]}),
    .mi({open_n23434,\t/memstraddress [21]}),
    .sr(rst_pad),
    .q({open_n23440,\t/memstraddress [21]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b22  (
    .a({_al_u2852_o,_al_u2852_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [22],\t/a/ID_memstraddr [22]}),
    .mi({open_n23452,\t/memstraddress [22]}),
    .sr(rst_pad),
    .q({open_n23458,\t/memstraddress [22]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b23  (
    .a({_al_u2849_o,_al_u2849_o}),
    .b({\t/a/instr/n12 [23],\t/a/instr/n12 [23]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2850_o,_al_u2850_o}),
    .mi({open_n23470,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23476,\t/memstraddress [23]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b24  (
    .a({_al_u2846_o,_al_u2846_o}),
    .b({\t/a/instr/n12 [24],\t/a/instr/n12 [24]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2847_o,_al_u2847_o}),
    .mi({open_n23488,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23494,\t/memstraddress [24]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b25  (
    .a({_al_u2843_o,_al_u2843_o}),
    .b({\t/a/instr/n12 [25],\t/a/instr/n12 [25]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2844_o,_al_u2844_o}),
    .mi({open_n23506,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23512,\t/memstraddress [25]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b26  (
    .a({_al_u2840_o,_al_u2840_o}),
    .b({\t/a/instr/n12 [26],\t/a/instr/n12 [26]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2841_o,_al_u2841_o}),
    .mi({open_n23524,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23530,\t/memstraddress [26]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b27  (
    .a({_al_u2838_o,_al_u2838_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [27],\t/a/ID_memstraddr [27]}),
    .mi({open_n23542,\t/memstraddress [27]}),
    .sr(rst_pad),
    .q({open_n23548,\t/memstraddress [27]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b28  (
    .a({_al_u2836_o,_al_u2836_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [28],\t/a/ID_memstraddr [28]}),
    .mi({open_n23560,\t/memstraddress [28]}),
    .sr(rst_pad),
    .q({open_n23566,\t/memstraddress [28]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b29  (
    .a({_al_u2833_o,_al_u2833_o}),
    .b({\t/a/instr/n12 [29],\t/a/instr/n12 [29]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2834_o,_al_u2834_o}),
    .mi({open_n23578,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23584,\t/memstraddress [29]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b3  (
    .a({_al_u2831_o,_al_u2831_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [3],\t/a/ID_memstraddr [3]}),
    .mi({open_n23596,\t/memstraddress [3]}),
    .sr(rst_pad),
    .q({open_n23602,\t/memstraddress [3]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b30  (
    .a({_al_u2828_o,_al_u2828_o}),
    .b({\t/a/instr/n12 [30],\t/a/instr/n12 [30]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2829_o,_al_u2829_o}),
    .mi({open_n23614,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23620,\t/memstraddress [30]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b31  (
    .a({_al_u2826_o,_al_u2826_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [31],\t/a/ID_memstraddr [31]}),
    .mi({open_n23632,\t/memstraddress [31]}),
    .sr(rst_pad),
    .q({open_n23638,\t/memstraddress [31]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b4  (
    .a({_al_u2824_o,_al_u2824_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [4],\t/a/ID_memstraddr [4]}),
    .mi({open_n23650,\t/memstraddress [4]}),
    .sr(rst_pad),
    .q({open_n23656,\t/memstraddress [4]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b5  (
    .a({_al_u2821_o,_al_u2821_o}),
    .b({\t/a/instr/n12 [5],\t/a/instr/n12 [5]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2822_o,_al_u2822_o}),
    .mi({open_n23668,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23674,\t/memstraddress [5]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b6  (
    .a({_al_u2819_o,_al_u2819_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [6],\t/a/ID_memstraddr [6]}),
    .mi({open_n23686,\t/memstraddress [6]}),
    .sr(rst_pad),
    .q({open_n23692,\t/memstraddress [6]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*~(D)*~(C)+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*~(C)+~((0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B))*D*C+(0*~(A)*~(B)+0*A*~(B)+~(0)*A*B+0*A*B)*D*C)"),
    //.LUT1("((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*~(D)*~(C)+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*~(C)+~((1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B))*D*C+(1*~(A)*~(B)+1*A*~(B)+~(1)*A*B+1*A*B)*D*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100000001000),
    .INIT_LUT1(16'b1111101100001011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b7  (
    .a({_al_u2817_o,_al_u2817_o}),
    .b({_al_u2807_o,_al_u2807_o}),
    .c({\t/a/condition/n0_lutinv ,\t/a/condition/n0_lutinv }),
    .clk(clock_pad),
    .d({\t/a/ID_memstraddr [7],\t/a/ID_memstraddr [7]}),
    .mi({open_n23704,\t/memstraddress [7]}),
    .sr(rst_pad),
    .q({open_n23710,\t/memstraddress [7]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b8  (
    .a({_al_u2814_o,_al_u2814_o}),
    .b({\t/a/instr/n12 [8],\t/a/instr/n12 [8]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2815_o,_al_u2815_o}),
    .mi({open_n23722,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23728,\t/memstraddress [8]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("(D*~(C*~A*~(~0*B)))"),
    //.LUT1("(D*~(C*~A*~(~1*B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111100000000),
    .INIT_LUT1(16'b1010111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/instr/reg0_b9  (
    .a({_al_u2811_o,_al_u2811_o}),
    .b({\t/a/instr/n12 [9],\t/a/instr/n12 [9]}),
    .c({_al_u2808_o,_al_u2808_o}),
    .clk(clock_pad),
    .d({_al_u2812_o,_al_u2812_o}),
    .mi({open_n23740,_al_u2109_o}),
    .sr(rst_pad),
    .q({open_n23746,\t/memstraddress [9]}));  // PC.v(60)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~((0*~C))*~(B)+D*(0*~C)*~(B)+~(D)*(0*~C)*B+D*(0*~C)*B))"),
    //.LUT1("~(~A*~(D*~((1*~C))*~(B)+D*(1*~C)*~(B)+~(D)*(1*~C)*B+D*(1*~C)*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1011111110101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b10  (
    .a({_al_u1902_o,_al_u1902_o}),
    .b({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .c({_al_u1903_o,_al_u1903_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [10],\t/a/MEM_aludat [10]}),
    .mi({open_n23758,i_data[10]}),
    .sr(rst_pad),
    .q({open_n23764,\t/a/reg_writedat [10]}));  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~B*~A*~(D*~C))"),
    //.LUT1("~(~A*~(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1110111111101110),
    .INIT_LUT1(16'b1111101111101010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b11|t/a/mem_wb/reg0_b9  (
    .a({_al_u1902_o,_al_u1902_o}),
    .b({\t/busarbitration/mux5_b0_sel_is_3_o ,_al_u1904_o}),
    .c({_al_u1940_o,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [11],\t/a/MEM_aludat [9]}),
    .sr(rst_pad),
    .q({\t/a/reg_writedat [11],\t/a/reg_writedat [9]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~((0*~C))*~(B)+D*(0*~C)*~(B)+~(D)*(0*~C)*B+D*(0*~C)*B))"),
    //.LUT1("~(~A*~(D*~((1*~C))*~(B)+D*(1*~C)*~(B)+~(D)*(1*~C)*B+D*(1*~C)*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1011111110101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b12  (
    .a({_al_u1902_o,_al_u1902_o}),
    .b({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .c({_al_u1903_o,_al_u1903_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [12],\t/a/MEM_aludat [12]}),
    .mi({open_n23794,i_data[12]}),
    .sr(rst_pad),
    .q({open_n23800,\t/a/reg_writedat [12]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~((0*~C))*~(B)+D*(0*~C)*~(B)+~(D)*(0*~C)*B+D*(0*~C)*B))"),
    //.LUT1("~(~A*~(D*~((1*~C))*~(B)+D*(1*~C)*~(B)+~(D)*(1*~C)*B+D*(1*~C)*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1011111110101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b13  (
    .a({_al_u1902_o,_al_u1902_o}),
    .b({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .c({_al_u1903_o,_al_u1903_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [13],\t/a/MEM_aludat [13]}),
    .mi({open_n23812,i_data[13]}),
    .sr(rst_pad),
    .q({open_n23818,\t/a/reg_writedat [13]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~((0*~C))*~(B)+D*(0*~C)*~(B)+~(D)*(0*~C)*B+D*(0*~C)*B))"),
    //.LUT1("~(~A*~(D*~((1*~C))*~(B)+D*(1*~C)*~(B)+~(D)*(1*~C)*B+D*(1*~C)*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101110101010),
    .INIT_LUT1(16'b1011111110101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b14  (
    .a({_al_u1902_o,_al_u1902_o}),
    .b({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .c({_al_u1903_o,_al_u1903_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [14],\t/a/MEM_aludat [14]}),
    .mi({open_n23830,i_data[14]}),
    .sr(rst_pad),
    .q({open_n23836,\t/a/reg_writedat [14]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b16  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [16],\t/a/MEM_aludat [16]}),
    .mi({open_n23848,i_data[16]}),
    .sr(rst_pad),
    .q({open_n23854,\t/a/reg_writedat [16]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b17  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [17],\t/a/MEM_aludat [17]}),
    .mi({open_n23866,i_data[17]}),
    .sr(rst_pad),
    .q({open_n23872,\t/a/reg_writedat [17]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b18  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [18],\t/a/MEM_aludat [18]}),
    .mi({open_n23884,i_data[18]}),
    .sr(rst_pad),
    .q({open_n23890,\t/a/reg_writedat [18]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b19  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [19],\t/a/MEM_aludat [19]}),
    .mi({open_n23902,i_data[19]}),
    .sr(rst_pad),
    .q({open_n23908,\t/a/reg_writedat [19]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b20  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [20],\t/a/MEM_aludat [20]}),
    .mi({open_n23920,i_data[20]}),
    .sr(rst_pad),
    .q({open_n23926,\t/a/reg_writedat [20]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b21  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [21],\t/a/MEM_aludat [21]}),
    .mi({open_n23938,i_data[21]}),
    .sr(rst_pad),
    .q({open_n23944,\t/a/reg_writedat [21]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b22  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [22],\t/a/MEM_aludat [22]}),
    .mi({open_n23956,i_data[22]}),
    .sr(rst_pad),
    .q({open_n23962,\t/a/reg_writedat [22]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b23  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [23],\t/a/MEM_aludat [23]}),
    .mi({open_n23974,i_data[23]}),
    .sr(rst_pad),
    .q({open_n23980,\t/a/reg_writedat [23]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b24  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [24],\t/a/MEM_aludat [24]}),
    .mi({open_n23992,i_data[24]}),
    .sr(rst_pad),
    .q({open_n23998,\t/a/reg_writedat [24]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b25  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [25],\t/a/MEM_aludat [25]}),
    .mi({open_n24010,i_data[25]}),
    .sr(rst_pad),
    .q({open_n24016,\t/a/reg_writedat [25]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b26  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [26],\t/a/MEM_aludat [26]}),
    .mi({open_n24028,i_data[26]}),
    .sr(rst_pad),
    .q({open_n24034,\t/a/reg_writedat [26]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b27  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [27],\t/a/MEM_aludat [27]}),
    .mi({open_n24046,i_data[27]}),
    .sr(rst_pad),
    .q({open_n24052,\t/a/reg_writedat [27]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b28  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [28],\t/a/MEM_aludat [28]}),
    .mi({open_n24064,i_data[28]}),
    .sr(rst_pad),
    .q({open_n24070,\t/a/reg_writedat [28]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b29  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [29],\t/a/MEM_aludat [29]}),
    .mi({open_n24082,i_data[29]}),
    .sr(rst_pad),
    .q({open_n24088,\t/a/reg_writedat [29]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b30  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [30],\t/a/MEM_aludat [30]}),
    .mi({open_n24100,i_data[30]}),
    .sr(rst_pad),
    .q({open_n24106,\t/a/reg_writedat [30]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(~A*~(D*~C)*~(0*B))"),
    //.LUT1("~(~A*~(D*~C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111110101010),
    .INIT_LUT1(16'b1110111111101110),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg0_b31  (
    .a({_al_u1917_o,_al_u1917_o}),
    .b({_al_u1918_o,_al_u1918_o}),
    .c({\t/busarbitration/mux5_b0_sel_is_3_o ,\t/busarbitration/mux5_b0_sel_is_3_o }),
    .clk(clock_pad),
    .d({\t/a/MEM_aludat [31],\t/a/MEM_aludat [31]}),
    .mi({open_n24118,i_data[31]}),
    .sr(rst_pad),
    .q({open_n24124,\t/a/reg_writedat [31]}));  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("(~D)"),
    //.LUT1("(~C*B*D)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011111111),
    .INIT_LUT1(16'b0000110000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \t/a/mem_wb/reg1_b1|t/a/mem_wb/reg1_b0  (
    .b({\t/a/MEM_op [1],open_n24127}),
    .c({\t/a/MEM_op [2],open_n24128}),
    .ce(\t/a/ex_mem/n0 ),
    .clk(clock_pad),
    .d({\t/a/MEM_op [0],rst_pad}),
    .mi(\t/a/MEM_op [1:0]),
    .f({_al_u251_o,\t/a/ex_mem/n0 }),
    .q(\t/a/WB_op [1:0]));  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~D)"),
    //.LUTF1("(D*~C*~B*~A)"),
    //.LUTG0("(~C*~D)"),
    //.LUTG1("(D*~C*~B*~A)"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001111),
    .INIT_LUTF1(16'b0000000100000000),
    .INIT_LUTG0(16'b0000000000001111),
    .INIT_LUTG1(16'b0000000100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \t/a/mem_wb/reg1_b2|t/a/mem_wb/reg1_b3  (
    .a({\t/a/WB_op [2],open_n24143}),
    .b({\t/a/WB_op [3],open_n24144}),
    .c({\t/a/WB_op [4],\t/a/MEM_op [4]}),
    .ce(\t/a/ex_mem/n0 ),
    .clk(clock_pad),
    .d({\t/a/WB_op [5],\t/a/MEM_op [3]}),
    .mi({\t/a/MEM_op [2],\t/a/MEM_op [3]}),
    .f({_al_u1793_o,_al_u252_o}),
    .q({\t/a/WB_op [2],\t/a/WB_op [3]}));  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \t/a/mem_wb/reg1_b4  (
    .ce(\t/a/ex_mem/n0 ),
    .clk(clock_pad),
    .mi({open_n24174,\t/a/MEM_op [4]}),
    .q({open_n24192,\t/a/WB_op [4]}));  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  // flow_line_reg.v(234)
  EG_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/reg2_b2|t/a/mem_wb/reg2_b0  (
    .a({_al_u1968_o,_al_u1967_o}),
    .b({_al_u1969_o,\t/a/MEM_rd [0]}),
    .c({_al_u1970_o,\t/a/MEM_rd [1]}),
    .clk(clock_pad),
    .d({\t/a/MEM_rd [2],\t/a/EX_rs2 [0]}),
    .e(\t/a/EX_rs2 [2:1]),
    .mi({\t/a/MEM_rd [2],\t/a/MEM_rd [0]}),
    .sr(rst_pad),
    .f({\t/a/n24_lutinv ,_al_u1968_o}),
    .q({\t/a/WB_rd [2],\t/a/WB_rd [0]}));  // flow_line_reg.v(234)
  EG_PHY_MSLICE #(
    //.LUT0("~(C*((~0*B)*~(A)*~(D)+(~0*B)*A*~(D)+~((~0*B))*A*D+(~0*B)*A*D))"),
    //.LUT1("~(C*((~1*B)*~(A)*~(D)+(~1*B)*A*~(D)+~((~1*B))*A*D+(~1*B)*A*D))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101111100111111),
    .INIT_LUT1(16'b0101111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/mem_wb/regwritecs_reg  (
    .a({_al_u251_o,_al_u251_o}),
    .b({_al_u290_o,_al_u290_o}),
    .c({_al_u252_o,_al_u252_o}),
    .clk(clock_pad),
    .d({\t/a/MEM_op [5],\t/a/MEM_op [5]}),
    .mi({open_n24220,\t/a/MEM_op [6]}),
    .sr(rst_pad),
    .q({open_n24226,\t/a/WB_regwritecs }));  // flow_line_reg.v(234)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b0|t/a/regfile/reg0_b9  (
    .a({open_n24227,\t/a/ID_rs2 [0]}),
    .b({open_n24228,\t/a/ID_rs2 [1]}),
    .c({\t/a/WB_regwritecs ,\t/a/regfile/regfile$1$ [9]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/n46 [0],\t/a/regfile/regfile$0$ [9]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [9]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b0_sel_is_3_o ,_al_u1052_o}),
    .q({\t/a/regfile/regfile$0$ [0],\t/a/regfile/regfile$0$ [9]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b1000|t/a/regfile/reg0_b999  (
    .a({_al_u256_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$30$ [7]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$31$ [7]}),
    .mi(\t/a/reg_writedat [8:7]),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b1000_sel_is_3_o ,_al_u1107_o}),
    .q(\t/a/regfile/regfile$31$ [8:7]));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0101000101000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0101000101000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b1001|t/a/regfile/reg0_b996  (
    .a({_al_u2614_o,\t/a/ID_rs2 [0]}),
    .b({_al_u2616_o,\t/a/ID_rs2 [1]}),
    .c({\t/a/MEM_aludat [9],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [9],\t/a/regfile/regfile$30$ [4]}),
    .e({open_n24257,\t/a/regfile/regfile$31$ [4]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u2718_o,_al_u1170_o}),
    .q({\t/a/regfile/regfile$31$ [9],\t/a/regfile/regfile$31$ [4]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b1002|t/a/regfile/reg0_b995  (
    .a({_al_u2606_o,\t/a/ID_rs2 [0]}),
    .b({_al_u2610_o,\t/a/ID_rs2 [1]}),
    .c({\t/a/MEM_aludat [10],\t/a/regfile/regfile$30$ [3]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [10],\t/a/regfile/regfile$31$ [3]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u2711_o,_al_u1177_o}),
    .q({\t/a/regfile/regfile$31$ [10],\t/a/regfile/regfile$31$ [3]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b101|t/a/regfile/reg0_b99  (
    .a({_al_u2614_o,\t/a/ID_rs2 [0]}),
    .b({_al_u2616_o,\t/a/ID_rs2 [1]}),
    .c({\t/a/MEM_aludat [5],\t/a/regfile/regfile$2$ [3]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [5],\t/a/regfile/regfile$3$ [3]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u2740_o,_al_u1189_o}),
    .q({\t/a/regfile/regfile$3$ [5],\t/a/regfile/regfile$3$ [3]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b102|t/a/regfile/reg0_b98  (
    .a({_al_u2614_o,\t/a/ID_rs2 [0]}),
    .b({_al_u2616_o,\t/a/ID_rs2 [1]}),
    .c({\t/a/MEM_aludat [6],\t/a/regfile/regfile$2$ [2]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [6],\t/a/regfile/regfile$3$ [2]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [2]}),
    .sr(rst_pad),
    .f({_al_u2733_o,_al_u1242_o}),
    .q({\t/a/regfile/regfile$3$ [6],\t/a/regfile/regfile$3$ [2]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b103|t/a/regfile/reg0_b97  (
    .a({_al_u2614_o,\t/a/ID_rs2 [0]}),
    .b({_al_u2616_o,\t/a/ID_rs2 [1]}),
    .c({\t/a/MEM_aludat [7],\t/a/regfile/regfile$2$ [1]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [7],\t/a/regfile/regfile$3$ [1]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [1]}),
    .sr(rst_pad),
    .f({_al_u2726_o,_al_u1473_o}),
    .q({\t/a/regfile/regfile$3$ [7],\t/a/regfile/regfile$3$ [1]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b107|t/a/regfile/reg0_b126  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/MEM_aludat [11],\t/a/MEM_aludat [30]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [11],\t/a/reg_writedat [30]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u2703_o,_al_u2619_o}),
    .q({\t/a/regfile/regfile$3$ [11],\t/a/regfile/regfile$3$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b108|t/a/regfile/reg0_b125  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/MEM_aludat [12],\t/a/MEM_aludat [29]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [12],\t/a/reg_writedat [29]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u2699_o,_al_u2623_o}),
    .q({\t/a/regfile/regfile$3$ [12],\t/a/regfile/regfile$3$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b109|t/a/regfile/reg0_b122  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/MEM_aludat [13],\t/a/MEM_aludat [26]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [13],\t/a/reg_writedat [26]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u2695_o,_al_u2635_o}),
    .q({\t/a/regfile/regfile$3$ [13],\t/a/regfile/regfile$3$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b10|t/a/regfile/reg0_b8  (
    .a({_al_u2614_o,\t/a/ID_rs2 [0]}),
    .b({_al_u2616_o,\t/a/ID_rs2 [1]}),
    .c({\t/a/MEM_aludat [10],\t/a/regfile/regfile$1$ [8]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [10],\t/a/regfile/regfile$0$ [8]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [8]}),
    .sr(rst_pad),
    .f({_al_u2714_o,_al_u1083_o}),
    .q({\t/a/regfile/regfile$0$ [10],\t/a/regfile/regfile$0$ [8]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b110|t/a/regfile/reg0_b121  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/MEM_aludat [14],\t/a/MEM_aludat [25]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [14],\t/a/reg_writedat [25]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u2689_o,_al_u2639_o}),
    .q({\t/a/regfile/regfile$3$ [14],\t/a/regfile/regfile$3$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b111|t/a/regfile/reg0_b118  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/MEM_aludat [15],\t/a/MEM_aludat [22]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [15],\t/a/reg_writedat [22]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u2681_o,_al_u2651_o}),
    .q({\t/a/regfile/regfile$3$ [15],\t/a/regfile/regfile$3$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b112|t/a/regfile/reg0_b117  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/MEM_aludat [16],\t/a/MEM_aludat [21]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [16],\t/a/reg_writedat [21]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u2675_o,_al_u2655_o}),
    .q({\t/a/regfile/regfile$3$ [16],\t/a/regfile/regfile$3$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000101000000),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b113|t/a/regfile/reg0_b114  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({_al_u2610_o,_al_u2610_o}),
    .c({\t/a/MEM_aludat [17],\t/a/MEM_aludat [18]}),
    .ce(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [17],\t/a/reg_writedat [18]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u2671_o,_al_u2667_o}),
    .q({\t/a/regfile/regfile$3$ [17],\t/a/regfile/regfile$3$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b11|t/a/regfile/reg0_b7  (
    .a({_al_u2066_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/alu_B_select [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/aluin/n10_lutinv ,\t/a/regfile/regfile$1$ [7]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [11],\t/a/regfile/regfile$0$ [7]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [7]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b11/B9 ,_al_u1094_o}),
    .q({\t/a/regfile/regfile$0$ [11],\t/a/regfile/regfile$0$ [7]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b12|t/a/regfile/reg0_b6  (
    .a({_al_u2063_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/alu_B_select [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/aluin/n10_lutinv ,\t/a/regfile/regfile$1$ [6]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [12],\t/a/regfile/regfile$0$ [6]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b12/B9 ,_al_u1115_o}),
    .q({\t/a/regfile/regfile$0$ [12],\t/a/regfile/regfile$0$ [6]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b137|t/a/regfile/reg0_b145  (
    .a({_al_u1979_o,_al_u2048_o}),
    .b({\t/a/alu_B_select [1],\t/a/alu_B_select [1]}),
    .c({\t/a/aluin/n10_lutinv ,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [9],\t/a/reg_writedat [17]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b9/B9 ,\t/a/aluin/sel1_b17/B9 }),
    .q({\t/a/regfile/regfile$4$ [9],\t/a/regfile/regfile$4$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b13|t/a/regfile/reg0_b5  (
    .a({_al_u2060_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/alu_B_select [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/aluin/n10_lutinv ,\t/a/regfile/regfile$1$ [5]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [13],\t/a/regfile/regfile$0$ [5]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b13/B9 ,_al_u1136_o}),
    .q({\t/a/regfile/regfile$0$ [13],\t/a/regfile/regfile$0$ [5]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(C*~A*~(~D*B))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101000000010000),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b143|t/a/regfile/reg0_b144  (
    .a({_al_u2054_o,_al_u2051_o}),
    .b({\t/a/alu_B_select [1],\t/a/alu_B_select [1]}),
    .c({\t/a/aluin/n10_lutinv ,\t/a/aluin/n10_lutinv }),
    .ce(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b15/B9 ,\t/a/aluin/sel1_b16/B9 }),
    .q({\t/a/regfile/regfile$4$ [15],\t/a/regfile/regfile$4$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000010011),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b14|t/a/regfile/reg0_b4  (
    .a({_al_u2057_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/alu_B_select [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/aluin/n10_lutinv ,\t/a/regfile/regfile$1$ [4]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [14],\t/a/regfile/regfile$0$ [4]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel1_b14/B9 ,_al_u1157_o}),
    .q({\t/a/regfile/regfile$0$ [14],\t/a/regfile/regfile$0$ [4]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b15|t/a/regfile/reg0_b31  (
    .a({_al_u1877_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$0$ [31]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [15],\t/a/regfile/regfile$1$ [31]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b15/B0 ,_al_u493_o}),
    .q({\t/a/regfile/regfile$0$ [15],\t/a/regfile/regfile$0$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b162|t/a/regfile/reg0_b177  (
    .a({_al_u2606_o,\t/a/ID_rs1 [0]}),
    .b({_al_u2610_o,\t/a/ID_rs1 [1]}),
    .c({\t/a/MEM_aludat [2],\t/a/regfile/regfile$4$ [17]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [2],\t/a/regfile/regfile$5$ [17]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u2754_o,_al_u817_o}),
    .q({\t/a/regfile/regfile$5$ [2],\t/a/regfile/regfile$5$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b163|t/a/regfile/reg0_b176  (
    .a({_al_u2606_o,\t/a/ID_rs1 [0]}),
    .b({_al_u2610_o,\t/a/ID_rs1 [1]}),
    .c({\t/a/MEM_aludat [3],\t/a/regfile/regfile$4$ [16]}),
    .ce(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [3],\t/a/regfile/regfile$5$ [16]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u2749_o,_al_u848_o}),
    .q({\t/a/regfile/regfile$5$ [3],\t/a/regfile/regfile$5$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b16|t/a/regfile/reg0_b30  (
    .a({_al_u1874_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$0$ [30]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [16],\t/a/regfile/regfile$1$ [30]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b16/B0 ,_al_u504_o}),
    .q({\t/a/regfile/regfile$0$ [16],\t/a/regfile/regfile$0$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b17|t/a/regfile/reg0_b3  (
    .a({_al_u1871_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$0$ [3]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [17],\t/a/regfile/regfile$1$ [3]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b17/B0 ,_al_u462_o}),
    .q({\t/a/regfile/regfile$0$ [17],\t/a/regfile/regfile$0$ [3]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b18|t/a/regfile/reg0_b29  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$0$ [18],\t/a/regfile/regfile$0$ [29]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [18],\t/a/regfile/regfile$1$ [29]}),
    .mi({\t/a/reg_writedat [18],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u808_o,_al_u556_o}),
    .q({\t/a/regfile/regfile$0$ [18],\t/a/regfile/regfile$0$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b193|t/a/regfile/reg0_b223  (
    .a({_al_u1895_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [31]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [1],\t/a/regfile/regfile$7$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b1/B0 ,_al_u492_o}),
    .q({\t/a/regfile/regfile$6$ [1],\t/a/regfile/regfile$6$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b197|t/a/regfile/reg0_b222  (
    .a({_al_u1817_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [30]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [5],\t/a/regfile/regfile$7$ [30]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b5/B0 ,_al_u503_o}),
    .q({\t/a/regfile/regfile$6$ [5],\t/a/regfile/regfile$6$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b198|t/a/regfile/reg0_b221  (
    .a({_al_u1814_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [29]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [6],\t/a/regfile/regfile$7$ [29]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b6/B0 ,_al_u555_o}),
    .q({\t/a/regfile/regfile$6$ [6],\t/a/regfile/regfile$6$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b199|t/a/regfile/reg0_b220  (
    .a({_al_u1811_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [28]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [7],\t/a/regfile/regfile$7$ [28]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b7/B0 ,_al_u566_o}),
    .q({\t/a/regfile/regfile$6$ [7],\t/a/regfile/regfile$6$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b19|t/a/regfile/reg0_b28  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$0$ [19],\t/a/regfile/regfile$0$ [28]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [19],\t/a/regfile/regfile$1$ [28]}),
    .mi({\t/a/reg_writedat [19],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u777_o,_al_u567_o}),
    .q({\t/a/regfile/regfile$0$ [19],\t/a/regfile/regfile$0$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101000101000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b1|t/a/regfile/reg0_b27  (
    .a({_al_u2614_o,\t/a/ID_rs1 [0]}),
    .b({_al_u2616_o,\t/a/ID_rs1 [1]}),
    .c({\t/a/MEM_aludat [1],\t/a/regfile/regfile$0$ [27]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [1],\t/a/regfile/regfile$1$ [27]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u2764_o,_al_u598_o}),
    .q({\t/a/regfile/regfile$0$ [1],\t/a/regfile/regfile$0$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b200|t/a/regfile/reg0_b219  (
    .a({_al_u1808_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [27]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [8],\t/a/regfile/regfile$7$ [27]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b8/B0 ,_al_u597_o}),
    .q({\t/a/regfile/regfile$6$ [8],\t/a/regfile/regfile$6$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b201|t/a/regfile/reg0_b218  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$6$ [9],\t/a/regfile/regfile$6$ [26]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [9],\t/a/regfile/regfile$7$ [26]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u345_o,_al_u608_o}),
    .q({\t/a/regfile/regfile$6$ [9],\t/a/regfile/regfile$6$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b202|t/a/regfile/reg0_b217  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$6$ [10],\t/a/regfile/regfile$6$ [25]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [10],\t/a/regfile/regfile$7$ [25]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u965_o,_al_u629_o}),
    .q({\t/a/regfile/regfile$6$ [10],\t/a/regfile/regfile$6$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b203|t/a/regfile/reg0_b216  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$6$ [11],\t/a/regfile/regfile$6$ [24]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [11],\t/a/regfile/regfile$7$ [24]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u954_o,_al_u650_o}),
    .q({\t/a/regfile/regfile$6$ [11],\t/a/regfile/regfile$6$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b204|t/a/regfile/reg0_b215  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$6$ [12],\t/a/regfile/regfile$6$ [23]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [12],\t/a/regfile/regfile$7$ [23]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u923_o,_al_u671_o}),
    .q({\t/a/regfile/regfile$6$ [12],\t/a/regfile/regfile$6$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b205|t/a/regfile/reg0_b214  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$6$ [13],\t/a/regfile/regfile$6$ [22]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [13],\t/a/regfile/regfile$7$ [22]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u912_o,_al_u702_o}),
    .q({\t/a/regfile/regfile$6$ [13],\t/a/regfile/regfile$6$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b206|t/a/regfile/reg0_b213  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$6$ [14],\t/a/regfile/regfile$6$ [21]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [14],\t/a/regfile/regfile$7$ [21]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u881_o,_al_u713_o}),
    .q({\t/a/regfile/regfile$6$ [14],\t/a/regfile/regfile$6$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b207|t/a/regfile/reg0_b212  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$6$ [15],\t/a/regfile/regfile$6$ [20]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [15],\t/a/regfile/regfile$7$ [20]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u860_o,_al_u744_o}),
    .q({\t/a/regfile/regfile$6$ [15],\t/a/regfile/regfile$6$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b208|t/a/regfile/reg0_b211  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$6$ [16],\t/a/regfile/regfile$6$ [19]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [16],\t/a/regfile/regfile$7$ [19]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u849_o,_al_u776_o}),
    .q({\t/a/regfile/regfile$6$ [16],\t/a/regfile/regfile$6$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b209|t/a/regfile/reg0_b210  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$6$ [17],\t/a/regfile/regfile$6$ [18]}),
    .ce(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [17],\t/a/regfile/regfile$7$ [18]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u818_o,_al_u807_o}),
    .q({\t/a/regfile/regfile$6$ [17],\t/a/regfile/regfile$6$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b20|t/a/regfile/reg0_b26  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$0$ [20],\t/a/regfile/regfile$0$ [26]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [20],\t/a/regfile/regfile$1$ [26]}),
    .mi({\t/a/reg_writedat [20],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u745_o,_al_u609_o}),
    .q({\t/a/regfile/regfile$0$ [20],\t/a/regfile/regfile$0$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b21|t/a/regfile/reg0_b25  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$0$ [21],\t/a/regfile/regfile$0$ [25]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [21],\t/a/regfile/regfile$1$ [25]}),
    .mi({\t/a/reg_writedat [21],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u714_o,_al_u630_o}),
    .q({\t/a/regfile/regfile$0$ [21],\t/a/regfile/regfile$0$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b225|t/a/regfile/reg0_b255  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [1],\t/a/regfile/regfile$6$ [31]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [1],\t/a/regfile/regfile$7$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u755_o,_al_u1198_o}),
    .q({\t/a/regfile/regfile$7$ [1],\t/a/regfile/regfile$7$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b226|t/a/regfile/reg0_b254  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [2],\t/a/regfile/regfile$6$ [30]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [2],\t/a/regfile/regfile$7$ [30]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u524_o,_al_u1229_o}),
    .q({\t/a/regfile/regfile$7$ [2],\t/a/regfile/regfile$7$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b227|t/a/regfile/reg0_b253  (
    .a({_al_u1829_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [29]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [3],\t/a/regfile/regfile$7$ [29]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b3/B0 ,_al_u1261_o}),
    .q({\t/a/regfile/regfile$7$ [3],\t/a/regfile/regfile$7$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b228|t/a/regfile/reg0_b252  (
    .a({_al_u1820_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$6$ [28]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [4],\t/a/regfile/regfile$7$ [28]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b4/B0 ,_al_u1292_o}),
    .q({\t/a/regfile/regfile$7$ [4],\t/a/regfile/regfile$7$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b229|t/a/regfile/reg0_b251  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [5],\t/a/regfile/regfile$6$ [27]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [5],\t/a/regfile/regfile$7$ [27]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u419_o,_al_u1303_o}),
    .q({\t/a/regfile/regfile$7$ [5],\t/a/regfile/regfile$7$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b22|t/a/regfile/reg0_b24  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$0$ [22],\t/a/regfile/regfile$0$ [24]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [22],\t/a/regfile/regfile$1$ [24]}),
    .mi({\t/a/reg_writedat [22],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u703_o,_al_u651_o}),
    .q({\t/a/regfile/regfile$0$ [22],\t/a/regfile/regfile$0$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b230|t/a/regfile/reg0_b250  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [6],\t/a/regfile/regfile$6$ [26]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [6],\t/a/regfile/regfile$7$ [26]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u398_o,_al_u1334_o}),
    .q({\t/a/regfile/regfile$7$ [6],\t/a/regfile/regfile$7$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b231|t/a/regfile/reg0_b249  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [7],\t/a/regfile/regfile$6$ [25]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [7],\t/a/regfile/regfile$7$ [25]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u387_o,_al_u1345_o}),
    .q({\t/a/regfile/regfile$7$ [7],\t/a/regfile/regfile$7$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b232|t/a/regfile/reg0_b248  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [8],\t/a/regfile/regfile$6$ [24]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [8],\t/a/regfile/regfile$7$ [24]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u356_o,_al_u1366_o}),
    .q({\t/a/regfile/regfile$7$ [8],\t/a/regfile/regfile$7$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b233|t/a/regfile/reg0_b247  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [9],\t/a/regfile/regfile$6$ [23]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [9],\t/a/regfile/regfile$7$ [23]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1051_o,_al_u1397_o}),
    .q({\t/a/regfile/regfile$7$ [9],\t/a/regfile/regfile$7$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b234|t/a/regfile/reg0_b246  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [10],\t/a/regfile/regfile$6$ [22]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [10],\t/a/regfile/regfile$7$ [22]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1691_o,_al_u1408_o}),
    .q({\t/a/regfile/regfile$7$ [10],\t/a/regfile/regfile$7$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b235|t/a/regfile/reg0_b245  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [11],\t/a/regfile/regfile$6$ [21]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [11],\t/a/regfile/regfile$7$ [21]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1660_o,_al_u1439_o}),
    .q({\t/a/regfile/regfile$7$ [11],\t/a/regfile/regfile$7$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b236|t/a/regfile/reg0_b244  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [12],\t/a/regfile/regfile$6$ [20]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [12],\t/a/regfile/regfile$7$ [20]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1649_o,_al_u1450_o}),
    .q({\t/a/regfile/regfile$7$ [12],\t/a/regfile/regfile$7$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b237|t/a/regfile/reg0_b243  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [13],\t/a/regfile/regfile$6$ [19]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [13],\t/a/regfile/regfile$7$ [19]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1618_o,_al_u1492_o}),
    .q({\t/a/regfile/regfile$7$ [13],\t/a/regfile/regfile$7$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b238|t/a/regfile/reg0_b242  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [14],\t/a/regfile/regfile$6$ [18]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [14],\t/a/regfile/regfile$7$ [18]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1597_o,_al_u1513_o}),
    .q({\t/a/regfile/regfile$7$ [14],\t/a/regfile/regfile$7$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b239|t/a/regfile/reg0_b241  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$6$ [15],\t/a/regfile/regfile$6$ [17]}),
    .ce(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$7$ [15],\t/a/regfile/regfile$7$ [17]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1586_o,_al_u1544_o}),
    .q({\t/a/regfile/regfile$7$ [15],\t/a/regfile/regfile$7$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b256|t/a/regfile/reg0_b287  (
    .a({_al_u254_o,_al_u498_o}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$8$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$9$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b256_sel_is_3_o ,_al_u499_o}),
    .q({\t/a/regfile/regfile$8$ [0],\t/a/regfile/regfile$8$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b257|t/a/regfile/reg0_b286  (
    .a({_al_u761_o,_al_u509_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [1],\t/a/regfile/regfile$8$ [30]}),
    .e({\t/a/regfile/regfile$9$ [1],\t/a/regfile/regfile$9$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u762_o,_al_u510_o}),
    .q({\t/a/regfile/regfile$8$ [1],\t/a/regfile/regfile$8$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b258|t/a/regfile/reg0_b285  (
    .a({_al_u530_o,_al_u561_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [2],\t/a/regfile/regfile$8$ [29]}),
    .e({\t/a/regfile/regfile$9$ [2],\t/a/regfile/regfile$9$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u531_o,_al_u562_o}),
    .q({\t/a/regfile/regfile$8$ [2],\t/a/regfile/regfile$8$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b259|t/a/regfile/reg0_b284  (
    .a({_al_u467_o,_al_u572_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [3],\t/a/regfile/regfile$8$ [28]}),
    .e({\t/a/regfile/regfile$9$ [3],\t/a/regfile/regfile$9$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u468_o,_al_u573_o}),
    .q({\t/a/regfile/regfile$8$ [3],\t/a/regfile/regfile$8$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b260|t/a/regfile/reg0_b283  (
    .a({_al_u456_o,_al_u603_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [4],\t/a/regfile/regfile$8$ [27]}),
    .e({\t/a/regfile/regfile$9$ [4],\t/a/regfile/regfile$9$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u457_o,_al_u604_o}),
    .q({\t/a/regfile/regfile$8$ [4],\t/a/regfile/regfile$8$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b261|t/a/regfile/reg0_b282  (
    .a({_al_u425_o,_al_u614_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [5],\t/a/regfile/regfile$8$ [26]}),
    .e({\t/a/regfile/regfile$9$ [5],\t/a/regfile/regfile$9$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u426_o,_al_u615_o}),
    .q({\t/a/regfile/regfile$8$ [5],\t/a/regfile/regfile$8$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b262|t/a/regfile/reg0_b281  (
    .a({_al_u404_o,_al_u635_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [6],\t/a/regfile/regfile$8$ [25]}),
    .e({\t/a/regfile/regfile$9$ [6],\t/a/regfile/regfile$9$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u405_o,_al_u636_o}),
    .q({\t/a/regfile/regfile$8$ [6],\t/a/regfile/regfile$8$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b263|t/a/regfile/reg0_b280  (
    .a({_al_u393_o,_al_u656_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [7],\t/a/regfile/regfile$8$ [24]}),
    .e({\t/a/regfile/regfile$9$ [7],\t/a/regfile/regfile$9$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u394_o,_al_u657_o}),
    .q({\t/a/regfile/regfile$8$ [7],\t/a/regfile/regfile$8$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b264|t/a/regfile/reg0_b279  (
    .a({_al_u362_o,_al_u677_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [8],\t/a/regfile/regfile$8$ [23]}),
    .e({\t/a/regfile/regfile$9$ [8],\t/a/regfile/regfile$9$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u363_o,_al_u678_o}),
    .q({\t/a/regfile/regfile$8$ [8],\t/a/regfile/regfile$8$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b265|t/a/regfile/reg0_b278  (
    .a({_al_u351_o,_al_u708_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [9],\t/a/regfile/regfile$8$ [22]}),
    .e({\t/a/regfile/regfile$9$ [9],\t/a/regfile/regfile$9$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u352_o,_al_u709_o}),
    .q({\t/a/regfile/regfile$8$ [9],\t/a/regfile/regfile$8$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b266|t/a/regfile/reg0_b277  (
    .a({_al_u971_o,_al_u719_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [10],\t/a/regfile/regfile$8$ [21]}),
    .e({\t/a/regfile/regfile$9$ [10],\t/a/regfile/regfile$9$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u972_o,_al_u720_o}),
    .q({\t/a/regfile/regfile$8$ [10],\t/a/regfile/regfile$8$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b267|t/a/regfile/reg0_b276  (
    .a({_al_u960_o,_al_u750_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [11],\t/a/regfile/regfile$8$ [20]}),
    .e({\t/a/regfile/regfile$9$ [11],\t/a/regfile/regfile$9$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u961_o,_al_u751_o}),
    .q({\t/a/regfile/regfile$8$ [11],\t/a/regfile/regfile$8$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b268|t/a/regfile/reg0_b275  (
    .a({_al_u929_o,_al_u782_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [12],\t/a/regfile/regfile$8$ [19]}),
    .e({\t/a/regfile/regfile$9$ [12],\t/a/regfile/regfile$9$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u930_o,_al_u783_o}),
    .q({\t/a/regfile/regfile$8$ [12],\t/a/regfile/regfile$8$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b269|t/a/regfile/reg0_b274  (
    .a({_al_u918_o,_al_u813_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [13],\t/a/regfile/regfile$8$ [18]}),
    .e({\t/a/regfile/regfile$9$ [13],\t/a/regfile/regfile$9$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u919_o,_al_u814_o}),
    .q({\t/a/regfile/regfile$8$ [13],\t/a/regfile/regfile$8$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b270|t/a/regfile/reg0_b273  (
    .a({_al_u887_o,_al_u824_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [14],\t/a/regfile/regfile$8$ [17]}),
    .e({\t/a/regfile/regfile$9$ [14],\t/a/regfile/regfile$9$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u888_o,_al_u825_o}),
    .q({\t/a/regfile/regfile$8$ [14],\t/a/regfile/regfile$8$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b271|t/a/regfile/reg0_b272  (
    .a({_al_u866_o,_al_u855_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [15],\t/a/regfile/regfile$8$ [16]}),
    .e({\t/a/regfile/regfile$9$ [15],\t/a/regfile/regfile$9$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u867_o,_al_u856_o}),
    .q({\t/a/regfile/regfile$8$ [15],\t/a/regfile/regfile$8$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*~D*~C*B*A)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*~D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b288|t/a/regfile/reg0_b319  (
    .a({_al_u254_o,_al_u1204_o}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$8$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$9$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b288_sel_is_3_o ,_al_u1205_o}),
    .q({\t/a/regfile/regfile$9$ [0],\t/a/regfile/regfile$9$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b289|t/a/regfile/reg0_b318  (
    .a({_al_u1477_o,_al_u1235_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [1],\t/a/regfile/regfile$8$ [30]}),
    .e({\t/a/regfile/regfile$9$ [1],\t/a/regfile/regfile$9$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1478_o,_al_u1236_o}),
    .q({\t/a/regfile/regfile$9$ [1],\t/a/regfile/regfile$9$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b290|t/a/regfile/reg0_b317  (
    .a({_al_u1246_o,_al_u1267_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [2],\t/a/regfile/regfile$8$ [29]}),
    .e({\t/a/regfile/regfile$9$ [2],\t/a/regfile/regfile$9$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1247_o,_al_u1268_o}),
    .q({\t/a/regfile/regfile$9$ [2],\t/a/regfile/regfile$9$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b291|t/a/regfile/reg0_b316  (
    .a({_al_u1193_o,_al_u1298_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [3],\t/a/regfile/regfile$8$ [28]}),
    .e({\t/a/regfile/regfile$9$ [3],\t/a/regfile/regfile$9$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1194_o,_al_u1299_o}),
    .q({\t/a/regfile/regfile$9$ [3],\t/a/regfile/regfile$9$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b292|t/a/regfile/reg0_b315  (
    .a({_al_u1162_o,_al_u1309_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [4],\t/a/regfile/regfile$8$ [27]}),
    .e({\t/a/regfile/regfile$9$ [4],\t/a/regfile/regfile$9$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1163_o,_al_u1310_o}),
    .q({\t/a/regfile/regfile$9$ [4],\t/a/regfile/regfile$9$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b293|t/a/regfile/reg0_b314  (
    .a({_al_u1141_o,_al_u1340_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [5],\t/a/regfile/regfile$8$ [26]}),
    .e({\t/a/regfile/regfile$9$ [5],\t/a/regfile/regfile$9$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1142_o,_al_u1341_o}),
    .q({\t/a/regfile/regfile$9$ [5],\t/a/regfile/regfile$9$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b294|t/a/regfile/reg0_b313  (
    .a({_al_u1120_o,_al_u1351_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [6],\t/a/regfile/regfile$8$ [25]}),
    .e({\t/a/regfile/regfile$9$ [6],\t/a/regfile/regfile$9$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1121_o,_al_u1352_o}),
    .q({\t/a/regfile/regfile$9$ [6],\t/a/regfile/regfile$9$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b295|t/a/regfile/reg0_b312  (
    .a({_al_u1099_o,_al_u1372_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [7],\t/a/regfile/regfile$8$ [24]}),
    .e({\t/a/regfile/regfile$9$ [7],\t/a/regfile/regfile$9$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1100_o,_al_u1373_o}),
    .q({\t/a/regfile/regfile$9$ [7],\t/a/regfile/regfile$9$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b296|t/a/regfile/reg0_b311  (
    .a({_al_u1088_o,_al_u1403_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [8],\t/a/regfile/regfile$8$ [23]}),
    .e({\t/a/regfile/regfile$9$ [8],\t/a/regfile/regfile$9$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1089_o,_al_u1404_o}),
    .q({\t/a/regfile/regfile$9$ [8],\t/a/regfile/regfile$9$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b297|t/a/regfile/reg0_b310  (
    .a({_al_u1057_o,_al_u1414_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [9],\t/a/regfile/regfile$8$ [22]}),
    .e({\t/a/regfile/regfile$9$ [9],\t/a/regfile/regfile$9$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1058_o,_al_u1415_o}),
    .q({\t/a/regfile/regfile$9$ [9],\t/a/regfile/regfile$9$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b298|t/a/regfile/reg0_b309  (
    .a({_al_u1697_o,_al_u1445_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [10],\t/a/regfile/regfile$8$ [21]}),
    .e({\t/a/regfile/regfile$9$ [10],\t/a/regfile/regfile$9$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1698_o,_al_u1446_o}),
    .q({\t/a/regfile/regfile$9$ [10],\t/a/regfile/regfile$9$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b299|t/a/regfile/reg0_b308  (
    .a({_al_u1666_o,_al_u1456_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [11],\t/a/regfile/regfile$8$ [20]}),
    .e({\t/a/regfile/regfile$9$ [11],\t/a/regfile/regfile$9$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1667_o,_al_u1457_o}),
    .q({\t/a/regfile/regfile$9$ [11],\t/a/regfile/regfile$9$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(C*~A*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0101000000010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b2|t/a/regfile/reg0_b23  (
    .a({_al_u1862_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/alu_A_select [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/aluin/n5_lutinv ,\t/a/regfile/regfile$0$ [23]}),
    .ce(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/reg_writedat [2],\t/a/regfile/regfile$1$ [23]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({\t/a/aluin/sel0_b2/B0 ,_al_u672_o}),
    .q({\t/a/regfile/regfile$0$ [2],\t/a/regfile/regfile$0$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b300|t/a/regfile/reg0_b307  (
    .a({_al_u1655_o,_al_u1498_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [12],\t/a/regfile/regfile$8$ [19]}),
    .e({\t/a/regfile/regfile$9$ [12],\t/a/regfile/regfile$9$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1656_o,_al_u1499_o}),
    .q({\t/a/regfile/regfile$9$ [12],\t/a/regfile/regfile$9$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b301|t/a/regfile/reg0_b306  (
    .a({_al_u1624_o,_al_u1519_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [13],\t/a/regfile/regfile$8$ [18]}),
    .e({\t/a/regfile/regfile$9$ [13],\t/a/regfile/regfile$9$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1625_o,_al_u1520_o}),
    .q({\t/a/regfile/regfile$9$ [13],\t/a/regfile/regfile$9$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b302|t/a/regfile/reg0_b305  (
    .a({_al_u1603_o,_al_u1550_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [14],\t/a/regfile/regfile$8$ [17]}),
    .e({\t/a/regfile/regfile$9$ [14],\t/a/regfile/regfile$9$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1604_o,_al_u1551_o}),
    .q({\t/a/regfile/regfile$9$ [14],\t/a/regfile/regfile$9$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b303|t/a/regfile/reg0_b304  (
    .a({_al_u1592_o,_al_u1561_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$8$ [15],\t/a/regfile/regfile$8$ [16]}),
    .e({\t/a/regfile/regfile$9$ [15],\t/a/regfile/regfile$9$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1593_o,_al_u1562_o}),
    .q({\t/a/regfile/regfile$9$ [15],\t/a/regfile/regfile$9$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*~D*C*~B*A)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*~D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b320|t/a/regfile/reg0_b351  (
    .a({_al_u254_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$10$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$11$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b320_sel_is_3_o ,_al_u498_o}),
    .q({\t/a/regfile/regfile$10$ [0],\t/a/regfile/regfile$10$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b321|t/a/regfile/reg0_b350  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [1],\t/a/regfile/regfile$10$ [30]}),
    .e({\t/a/regfile/regfile$11$ [1],\t/a/regfile/regfile$11$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u761_o,_al_u509_o}),
    .q({\t/a/regfile/regfile$10$ [1],\t/a/regfile/regfile$10$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b322|t/a/regfile/reg0_b349  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [2],\t/a/regfile/regfile$10$ [29]}),
    .e({\t/a/regfile/regfile$11$ [2],\t/a/regfile/regfile$11$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u530_o,_al_u561_o}),
    .q({\t/a/regfile/regfile$10$ [2],\t/a/regfile/regfile$10$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b323|t/a/regfile/reg0_b348  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [3],\t/a/regfile/regfile$10$ [28]}),
    .e({\t/a/regfile/regfile$11$ [3],\t/a/regfile/regfile$11$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u467_o,_al_u572_o}),
    .q({\t/a/regfile/regfile$10$ [3],\t/a/regfile/regfile$10$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b324|t/a/regfile/reg0_b347  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [4],\t/a/regfile/regfile$10$ [27]}),
    .e({\t/a/regfile/regfile$11$ [4],\t/a/regfile/regfile$11$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u456_o,_al_u603_o}),
    .q({\t/a/regfile/regfile$10$ [4],\t/a/regfile/regfile$10$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b325|t/a/regfile/reg0_b346  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [5],\t/a/regfile/regfile$10$ [26]}),
    .e({\t/a/regfile/regfile$11$ [5],\t/a/regfile/regfile$11$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u425_o,_al_u614_o}),
    .q({\t/a/regfile/regfile$10$ [5],\t/a/regfile/regfile$10$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b326|t/a/regfile/reg0_b345  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [6],\t/a/regfile/regfile$10$ [25]}),
    .e({\t/a/regfile/regfile$11$ [6],\t/a/regfile/regfile$11$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u404_o,_al_u635_o}),
    .q({\t/a/regfile/regfile$10$ [6],\t/a/regfile/regfile$10$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b327|t/a/regfile/reg0_b344  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [7],\t/a/regfile/regfile$10$ [24]}),
    .e({\t/a/regfile/regfile$11$ [7],\t/a/regfile/regfile$11$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u393_o,_al_u656_o}),
    .q({\t/a/regfile/regfile$10$ [7],\t/a/regfile/regfile$10$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b328|t/a/regfile/reg0_b343  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [8],\t/a/regfile/regfile$10$ [23]}),
    .e({\t/a/regfile/regfile$11$ [8],\t/a/regfile/regfile$11$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u362_o,_al_u677_o}),
    .q({\t/a/regfile/regfile$10$ [8],\t/a/regfile/regfile$10$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b329|t/a/regfile/reg0_b342  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [9],\t/a/regfile/regfile$10$ [22]}),
    .e({\t/a/regfile/regfile$11$ [9],\t/a/regfile/regfile$11$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u351_o,_al_u708_o}),
    .q({\t/a/regfile/regfile$10$ [9],\t/a/regfile/regfile$10$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b330|t/a/regfile/reg0_b341  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [10],\t/a/regfile/regfile$10$ [21]}),
    .e({\t/a/regfile/regfile$11$ [10],\t/a/regfile/regfile$11$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u971_o,_al_u719_o}),
    .q({\t/a/regfile/regfile$10$ [10],\t/a/regfile/regfile$10$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b331|t/a/regfile/reg0_b340  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [11],\t/a/regfile/regfile$10$ [20]}),
    .e({\t/a/regfile/regfile$11$ [11],\t/a/regfile/regfile$11$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u960_o,_al_u750_o}),
    .q({\t/a/regfile/regfile$10$ [11],\t/a/regfile/regfile$10$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b332|t/a/regfile/reg0_b339  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [12],\t/a/regfile/regfile$10$ [19]}),
    .e({\t/a/regfile/regfile$11$ [12],\t/a/regfile/regfile$11$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u929_o,_al_u782_o}),
    .q({\t/a/regfile/regfile$10$ [12],\t/a/regfile/regfile$10$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b333|t/a/regfile/reg0_b338  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [13],\t/a/regfile/regfile$10$ [18]}),
    .e({\t/a/regfile/regfile$11$ [13],\t/a/regfile/regfile$11$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u918_o,_al_u813_o}),
    .q({\t/a/regfile/regfile$10$ [13],\t/a/regfile/regfile$10$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b334|t/a/regfile/reg0_b337  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [14],\t/a/regfile/regfile$10$ [17]}),
    .e({\t/a/regfile/regfile$11$ [14],\t/a/regfile/regfile$11$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u887_o,_al_u824_o}),
    .q({\t/a/regfile/regfile$10$ [14],\t/a/regfile/regfile$10$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b335|t/a/regfile/reg0_b336  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [15],\t/a/regfile/regfile$10$ [16]}),
    .e({\t/a/regfile/regfile$11$ [15],\t/a/regfile/regfile$11$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u866_o,_al_u855_o}),
    .q({\t/a/regfile/regfile$10$ [15],\t/a/regfile/regfile$10$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b33|t/a/regfile/reg0_b63  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$0$ [1],\t/a/regfile/regfile$0$ [31]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [1],\t/a/regfile/regfile$1$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u756_o,_al_u1199_o}),
    .q({\t/a/regfile/regfile$1$ [1],\t/a/regfile/regfile$1$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b34|t/a/regfile/reg0_b62  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$0$ [2],\t/a/regfile/regfile$0$ [30]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [2],\t/a/regfile/regfile$1$ [30]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u525_o,_al_u1230_o}),
    .q({\t/a/regfile/regfile$1$ [2],\t/a/regfile/regfile$1$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*~D*C*B*A)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b352|t/a/regfile/reg0_b383  (
    .a({_al_u254_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$10$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$11$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b352_sel_is_3_o ,_al_u1204_o}),
    .q({\t/a/regfile/regfile$11$ [0],\t/a/regfile/regfile$11$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b353|t/a/regfile/reg0_b382  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [1],\t/a/regfile/regfile$10$ [30]}),
    .e({\t/a/regfile/regfile$11$ [1],\t/a/regfile/regfile$11$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1477_o,_al_u1235_o}),
    .q({\t/a/regfile/regfile$11$ [1],\t/a/regfile/regfile$11$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b354|t/a/regfile/reg0_b381  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [2],\t/a/regfile/regfile$10$ [29]}),
    .e({\t/a/regfile/regfile$11$ [2],\t/a/regfile/regfile$11$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1246_o,_al_u1267_o}),
    .q({\t/a/regfile/regfile$11$ [2],\t/a/regfile/regfile$11$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b355|t/a/regfile/reg0_b380  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [3],\t/a/regfile/regfile$10$ [28]}),
    .e({\t/a/regfile/regfile$11$ [3],\t/a/regfile/regfile$11$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1193_o,_al_u1298_o}),
    .q({\t/a/regfile/regfile$11$ [3],\t/a/regfile/regfile$11$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b356|t/a/regfile/reg0_b379  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [4],\t/a/regfile/regfile$10$ [27]}),
    .e({\t/a/regfile/regfile$11$ [4],\t/a/regfile/regfile$11$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1162_o,_al_u1309_o}),
    .q({\t/a/regfile/regfile$11$ [4],\t/a/regfile/regfile$11$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b357|t/a/regfile/reg0_b378  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [5],\t/a/regfile/regfile$10$ [26]}),
    .e({\t/a/regfile/regfile$11$ [5],\t/a/regfile/regfile$11$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1141_o,_al_u1340_o}),
    .q({\t/a/regfile/regfile$11$ [5],\t/a/regfile/regfile$11$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b358|t/a/regfile/reg0_b377  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [6],\t/a/regfile/regfile$10$ [25]}),
    .e({\t/a/regfile/regfile$11$ [6],\t/a/regfile/regfile$11$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1120_o,_al_u1351_o}),
    .q({\t/a/regfile/regfile$11$ [6],\t/a/regfile/regfile$11$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b359|t/a/regfile/reg0_b376  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [7],\t/a/regfile/regfile$10$ [24]}),
    .e({\t/a/regfile/regfile$11$ [7],\t/a/regfile/regfile$11$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1099_o,_al_u1372_o}),
    .q({\t/a/regfile/regfile$11$ [7],\t/a/regfile/regfile$11$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b35|t/a/regfile/reg0_b61  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$0$ [3],\t/a/regfile/regfile$0$ [29]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [3],\t/a/regfile/regfile$1$ [29]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1188_o,_al_u1262_o}),
    .q({\t/a/regfile/regfile$1$ [3],\t/a/regfile/regfile$1$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b360|t/a/regfile/reg0_b375  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [8],\t/a/regfile/regfile$10$ [23]}),
    .e({\t/a/regfile/regfile$11$ [8],\t/a/regfile/regfile$11$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1088_o,_al_u1403_o}),
    .q({\t/a/regfile/regfile$11$ [8],\t/a/regfile/regfile$11$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b361|t/a/regfile/reg0_b374  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [9],\t/a/regfile/regfile$10$ [22]}),
    .e({\t/a/regfile/regfile$11$ [9],\t/a/regfile/regfile$11$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1057_o,_al_u1414_o}),
    .q({\t/a/regfile/regfile$11$ [9],\t/a/regfile/regfile$11$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b362|t/a/regfile/reg0_b373  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [10],\t/a/regfile/regfile$10$ [21]}),
    .e({\t/a/regfile/regfile$11$ [10],\t/a/regfile/regfile$11$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1697_o,_al_u1445_o}),
    .q({\t/a/regfile/regfile$11$ [10],\t/a/regfile/regfile$11$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b363|t/a/regfile/reg0_b372  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [11],\t/a/regfile/regfile$10$ [20]}),
    .e({\t/a/regfile/regfile$11$ [11],\t/a/regfile/regfile$11$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1666_o,_al_u1456_o}),
    .q({\t/a/regfile/regfile$11$ [11],\t/a/regfile/regfile$11$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b364|t/a/regfile/reg0_b371  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [12],\t/a/regfile/regfile$10$ [19]}),
    .e({\t/a/regfile/regfile$11$ [12],\t/a/regfile/regfile$11$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1655_o,_al_u1498_o}),
    .q({\t/a/regfile/regfile$11$ [12],\t/a/regfile/regfile$11$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b365|t/a/regfile/reg0_b370  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [13],\t/a/regfile/regfile$10$ [18]}),
    .e({\t/a/regfile/regfile$11$ [13],\t/a/regfile/regfile$11$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1624_o,_al_u1519_o}),
    .q({\t/a/regfile/regfile$11$ [13],\t/a/regfile/regfile$11$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b366|t/a/regfile/reg0_b369  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [14],\t/a/regfile/regfile$10$ [17]}),
    .e({\t/a/regfile/regfile$11$ [14],\t/a/regfile/regfile$11$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1603_o,_al_u1550_o}),
    .q({\t/a/regfile/regfile$11$ [14],\t/a/regfile/regfile$11$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b367|t/a/regfile/reg0_b368  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$10$ [15],\t/a/regfile/regfile$10$ [16]}),
    .e({\t/a/regfile/regfile$11$ [15],\t/a/regfile/regfile$11$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1592_o,_al_u1561_o}),
    .q({\t/a/regfile/regfile$11$ [15],\t/a/regfile/regfile$11$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b36|t/a/regfile/reg0_b60  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$1$ [4],\t/a/regfile/regfile$0$ [28]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$0$ [4],\t/a/regfile/regfile$1$ [28]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u451_o,_al_u1293_o}),
    .q({\t/a/regfile/regfile$1$ [4],\t/a/regfile/regfile$1$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b37|t/a/regfile/reg0_b59  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$1$ [5],\t/a/regfile/regfile$0$ [27]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$0$ [5],\t/a/regfile/regfile$1$ [27]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u420_o,_al_u1304_o}),
    .q({\t/a/regfile/regfile$1$ [5],\t/a/regfile/regfile$1$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b38|t/a/regfile/reg0_b58  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$1$ [6],\t/a/regfile/regfile$0$ [26]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$0$ [6],\t/a/regfile/regfile$1$ [26]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u399_o,_al_u1335_o}),
    .q({\t/a/regfile/regfile$1$ [6],\t/a/regfile/regfile$1$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b39|t/a/regfile/reg0_b57  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$1$ [7],\t/a/regfile/regfile$0$ [25]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$0$ [7],\t/a/regfile/regfile$1$ [25]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u388_o,_al_u1346_o}),
    .q({\t/a/regfile/regfile$1$ [7],\t/a/regfile/regfile$1$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b40|t/a/regfile/reg0_b56  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$1$ [8],\t/a/regfile/regfile$0$ [24]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$0$ [8],\t/a/regfile/regfile$1$ [24]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u357_o,_al_u1367_o}),
    .q({\t/a/regfile/regfile$1$ [8],\t/a/regfile/regfile$1$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000001000010011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b41|t/a/regfile/reg0_b55  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$1$ [9],\t/a/regfile/regfile$0$ [23]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$0$ [9],\t/a/regfile/regfile$1$ [23]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u346_o,_al_u1398_o}),
    .q({\t/a/regfile/regfile$1$ [9],\t/a/regfile/regfile$1$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b42|t/a/regfile/reg0_b54  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$0$ [10],\t/a/regfile/regfile$0$ [22]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [10],\t/a/regfile/regfile$1$ [22]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u966_o,_al_u1409_o}),
    .q({\t/a/regfile/regfile$1$ [10],\t/a/regfile/regfile$1$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b43|t/a/regfile/reg0_b53  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$0$ [11],\t/a/regfile/regfile$0$ [21]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [11],\t/a/regfile/regfile$1$ [21]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u955_o,_al_u1440_o}),
    .q({\t/a/regfile/regfile$1$ [11],\t/a/regfile/regfile$1$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*D*C*~B*A)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b448|t/a/regfile/reg0_b479  (
    .a({_al_u254_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$14$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$15$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b448_sel_is_3_o ,_al_u496_o}),
    .q({\t/a/regfile/regfile$14$ [0],\t/a/regfile/regfile$14$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b449|t/a/regfile/reg0_b478  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [1],\t/a/regfile/regfile$14$ [30]}),
    .e({\t/a/regfile/regfile$15$ [1],\t/a/regfile/regfile$15$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u759_o,_al_u507_o}),
    .q({\t/a/regfile/regfile$14$ [1],\t/a/regfile/regfile$14$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b44|t/a/regfile/reg0_b52  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$0$ [12],\t/a/regfile/regfile$0$ [20]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [12],\t/a/regfile/regfile$1$ [20]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u924_o,_al_u1451_o}),
    .q({\t/a/regfile/regfile$1$ [12],\t/a/regfile/regfile$1$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b450|t/a/regfile/reg0_b477  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [2],\t/a/regfile/regfile$14$ [29]}),
    .e({\t/a/regfile/regfile$15$ [2],\t/a/regfile/regfile$15$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u528_o,_al_u559_o}),
    .q({\t/a/regfile/regfile$14$ [2],\t/a/regfile/regfile$14$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b451|t/a/regfile/reg0_b476  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [3],\t/a/regfile/regfile$14$ [28]}),
    .e({\t/a/regfile/regfile$15$ [3],\t/a/regfile/regfile$15$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u465_o,_al_u570_o}),
    .q({\t/a/regfile/regfile$14$ [3],\t/a/regfile/regfile$14$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b452|t/a/regfile/reg0_b475  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [4],\t/a/regfile/regfile$14$ [27]}),
    .e({\t/a/regfile/regfile$15$ [4],\t/a/regfile/regfile$15$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u454_o,_al_u601_o}),
    .q({\t/a/regfile/regfile$14$ [4],\t/a/regfile/regfile$14$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b453|t/a/regfile/reg0_b474  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [5],\t/a/regfile/regfile$14$ [26]}),
    .e({\t/a/regfile/regfile$15$ [5],\t/a/regfile/regfile$15$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u423_o,_al_u612_o}),
    .q({\t/a/regfile/regfile$14$ [5],\t/a/regfile/regfile$14$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b454|t/a/regfile/reg0_b473  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [6],\t/a/regfile/regfile$14$ [25]}),
    .e({\t/a/regfile/regfile$15$ [6],\t/a/regfile/regfile$15$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u402_o,_al_u633_o}),
    .q({\t/a/regfile/regfile$14$ [6],\t/a/regfile/regfile$14$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b455|t/a/regfile/reg0_b472  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [7],\t/a/regfile/regfile$14$ [24]}),
    .e({\t/a/regfile/regfile$15$ [7],\t/a/regfile/regfile$15$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u391_o,_al_u654_o}),
    .q({\t/a/regfile/regfile$14$ [7],\t/a/regfile/regfile$14$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b456|t/a/regfile/reg0_b471  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [8],\t/a/regfile/regfile$14$ [23]}),
    .e({\t/a/regfile/regfile$15$ [8],\t/a/regfile/regfile$15$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u360_o,_al_u675_o}),
    .q({\t/a/regfile/regfile$14$ [8],\t/a/regfile/regfile$14$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b457|t/a/regfile/reg0_b470  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [9],\t/a/regfile/regfile$14$ [22]}),
    .e({\t/a/regfile/regfile$15$ [9],\t/a/regfile/regfile$15$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u349_o,_al_u706_o}),
    .q({\t/a/regfile/regfile$14$ [9],\t/a/regfile/regfile$14$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b458|t/a/regfile/reg0_b469  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [10],\t/a/regfile/regfile$14$ [21]}),
    .e({\t/a/regfile/regfile$15$ [10],\t/a/regfile/regfile$15$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u969_o,_al_u717_o}),
    .q({\t/a/regfile/regfile$14$ [10],\t/a/regfile/regfile$14$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b459|t/a/regfile/reg0_b468  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [11],\t/a/regfile/regfile$14$ [20]}),
    .e({\t/a/regfile/regfile$15$ [11],\t/a/regfile/regfile$15$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u958_o,_al_u748_o}),
    .q({\t/a/regfile/regfile$14$ [11],\t/a/regfile/regfile$14$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b45|t/a/regfile/reg0_b51  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$0$ [13],\t/a/regfile/regfile$0$ [19]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [13],\t/a/regfile/regfile$1$ [19]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u913_o,_al_u1493_o}),
    .q({\t/a/regfile/regfile$1$ [13],\t/a/regfile/regfile$1$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b460|t/a/regfile/reg0_b467  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [12],\t/a/regfile/regfile$14$ [19]}),
    .e({\t/a/regfile/regfile$15$ [12],\t/a/regfile/regfile$15$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u927_o,_al_u780_o}),
    .q({\t/a/regfile/regfile$14$ [12],\t/a/regfile/regfile$14$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b461|t/a/regfile/reg0_b466  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [13],\t/a/regfile/regfile$14$ [18]}),
    .e({\t/a/regfile/regfile$15$ [13],\t/a/regfile/regfile$15$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u916_o,_al_u811_o}),
    .q({\t/a/regfile/regfile$14$ [13],\t/a/regfile/regfile$14$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b462|t/a/regfile/reg0_b465  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [14],\t/a/regfile/regfile$14$ [17]}),
    .e({\t/a/regfile/regfile$15$ [14],\t/a/regfile/regfile$15$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u885_o,_al_u822_o}),
    .q({\t/a/regfile/regfile$14$ [14],\t/a/regfile/regfile$14$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b463|t/a/regfile/reg0_b464  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [15],\t/a/regfile/regfile$14$ [16]}),
    .e({\t/a/regfile/regfile$15$ [15],\t/a/regfile/regfile$15$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u864_o,_al_u853_o}),
    .q({\t/a/regfile/regfile$14$ [15],\t/a/regfile/regfile$14$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b46|t/a/regfile/reg0_b50  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$0$ [14],\t/a/regfile/regfile$0$ [18]}),
    .ce(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$1$ [14],\t/a/regfile/regfile$1$ [18]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u882_o,_al_u1514_o}),
    .q({\t/a/regfile/regfile$1$ [14],\t/a/regfile/regfile$1$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b480|t/a/regfile/reg0_b511  (
    .a({_al_u254_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$14$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$15$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b480_sel_is_3_o ,_al_u1202_o}),
    .q({\t/a/regfile/regfile$15$ [0],\t/a/regfile/regfile$15$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b481|t/a/regfile/reg0_b510  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [1],\t/a/regfile/regfile$14$ [30]}),
    .e({\t/a/regfile/regfile$15$ [1],\t/a/regfile/regfile$15$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1475_o,_al_u1233_o}),
    .q({\t/a/regfile/regfile$15$ [1],\t/a/regfile/regfile$15$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b482|t/a/regfile/reg0_b509  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [2],\t/a/regfile/regfile$14$ [29]}),
    .e({\t/a/regfile/regfile$15$ [2],\t/a/regfile/regfile$15$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1244_o,_al_u1265_o}),
    .q({\t/a/regfile/regfile$15$ [2],\t/a/regfile/regfile$15$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b483|t/a/regfile/reg0_b508  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [3],\t/a/regfile/regfile$14$ [28]}),
    .e({\t/a/regfile/regfile$15$ [3],\t/a/regfile/regfile$15$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1191_o,_al_u1296_o}),
    .q({\t/a/regfile/regfile$15$ [3],\t/a/regfile/regfile$15$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b484|t/a/regfile/reg0_b507  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [4],\t/a/regfile/regfile$14$ [27]}),
    .e({\t/a/regfile/regfile$15$ [4],\t/a/regfile/regfile$15$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1160_o,_al_u1307_o}),
    .q({\t/a/regfile/regfile$15$ [4],\t/a/regfile/regfile$15$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b485|t/a/regfile/reg0_b506  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [5],\t/a/regfile/regfile$14$ [26]}),
    .e({\t/a/regfile/regfile$15$ [5],\t/a/regfile/regfile$15$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1139_o,_al_u1338_o}),
    .q({\t/a/regfile/regfile$15$ [5],\t/a/regfile/regfile$15$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b486|t/a/regfile/reg0_b505  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [6],\t/a/regfile/regfile$14$ [25]}),
    .e({\t/a/regfile/regfile$15$ [6],\t/a/regfile/regfile$15$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1118_o,_al_u1349_o}),
    .q({\t/a/regfile/regfile$15$ [6],\t/a/regfile/regfile$15$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b487|t/a/regfile/reg0_b504  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [7],\t/a/regfile/regfile$14$ [24]}),
    .e({\t/a/regfile/regfile$15$ [7],\t/a/regfile/regfile$15$ [24]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1097_o,_al_u1370_o}),
    .q({\t/a/regfile/regfile$15$ [7],\t/a/regfile/regfile$15$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b488|t/a/regfile/reg0_b503  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [8],\t/a/regfile/regfile$14$ [23]}),
    .e({\t/a/regfile/regfile$15$ [8],\t/a/regfile/regfile$15$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1086_o,_al_u1401_o}),
    .q({\t/a/regfile/regfile$15$ [8],\t/a/regfile/regfile$15$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b489|t/a/regfile/reg0_b502  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [9],\t/a/regfile/regfile$14$ [22]}),
    .e({\t/a/regfile/regfile$15$ [9],\t/a/regfile/regfile$15$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1055_o,_al_u1412_o}),
    .q({\t/a/regfile/regfile$15$ [9],\t/a/regfile/regfile$15$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b490|t/a/regfile/reg0_b501  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [10],\t/a/regfile/regfile$14$ [21]}),
    .e({\t/a/regfile/regfile$15$ [10],\t/a/regfile/regfile$15$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1695_o,_al_u1443_o}),
    .q({\t/a/regfile/regfile$15$ [10],\t/a/regfile/regfile$15$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b491|t/a/regfile/reg0_b500  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [11],\t/a/regfile/regfile$14$ [20]}),
    .e({\t/a/regfile/regfile$15$ [11],\t/a/regfile/regfile$15$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1664_o,_al_u1454_o}),
    .q({\t/a/regfile/regfile$15$ [11],\t/a/regfile/regfile$15$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b492|t/a/regfile/reg0_b499  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [12],\t/a/regfile/regfile$14$ [19]}),
    .e({\t/a/regfile/regfile$15$ [12],\t/a/regfile/regfile$15$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1653_o,_al_u1496_o}),
    .q({\t/a/regfile/regfile$15$ [12],\t/a/regfile/regfile$15$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b493|t/a/regfile/reg0_b498  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [13],\t/a/regfile/regfile$14$ [18]}),
    .e({\t/a/regfile/regfile$15$ [13],\t/a/regfile/regfile$15$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1622_o,_al_u1517_o}),
    .q({\t/a/regfile/regfile$15$ [13],\t/a/regfile/regfile$15$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b494|t/a/regfile/reg0_b497  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [14],\t/a/regfile/regfile$14$ [17]}),
    .e({\t/a/regfile/regfile$15$ [14],\t/a/regfile/regfile$15$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1601_o,_al_u1548_o}),
    .q({\t/a/regfile/regfile$15$ [14],\t/a/regfile/regfile$15$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b495|t/a/regfile/reg0_b496  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$14$ [15],\t/a/regfile/regfile$14$ [16]}),
    .e({\t/a/regfile/regfile$15$ [15],\t/a/regfile/regfile$15$ [16]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1590_o,_al_u1559_o}),
    .q({\t/a/regfile/regfile$15$ [15],\t/a/regfile/regfile$15$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b512|t/a/regfile/reg0_b543  (
    .a({_al_u256_o,_al_u488_o}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$16$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$17$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b512_sel_is_3_o ,_al_u489_o}),
    .q({\t/a/regfile/regfile$16$ [0],\t/a/regfile/regfile$16$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b513|t/a/regfile/reg0_b541  (
    .a({\t/a/ID_rs1 [0],_al_u551_o}),
    .b(\t/a/ID_rs1 [1:0]),
    .c({\t/a/regfile/regfile$16$ [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [1],\t/a/regfile/regfile$16$ [29]}),
    .e({open_n26677,\t/a/regfile/regfile$17$ [29]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u766_o,_al_u552_o}),
    .q({\t/a/regfile/regfile$16$ [1],\t/a/regfile/regfile$16$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b514|t/a/regfile/reg0_b539  (
    .a({\t/a/ID_rs1 [0],_al_u593_o}),
    .b(\t/a/ID_rs1 [1:0]),
    .c({\t/a/regfile/regfile$16$ [2],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [2],\t/a/regfile/regfile$16$ [27]}),
    .e({open_n26693,\t/a/regfile/regfile$17$ [27]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u535_o,_al_u594_o}),
    .q({\t/a/regfile/regfile$16$ [2],\t/a/regfile/regfile$16$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b515|t/a/regfile/reg0_b534  (
    .a({\t/a/ID_rs1 [0],_al_u698_o}),
    .b(\t/a/ID_rs1 [1:0]),
    .c({\t/a/regfile/regfile$16$ [3],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [3],\t/a/regfile/regfile$16$ [22]}),
    .e({open_n26709,\t/a/regfile/regfile$17$ [22]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u472_o,_al_u699_o}),
    .q({\t/a/regfile/regfile$16$ [3],\t/a/regfile/regfile$16$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b516|t/a/regfile/reg0_b532  (
    .a({_al_u446_o,_al_u740_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$16$ [4],\t/a/regfile/regfile$16$ [20]}),
    .e({\t/a/regfile/regfile$17$ [4],\t/a/regfile/regfile$17$ [20]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u447_o,_al_u741_o}),
    .q({\t/a/regfile/regfile$16$ [4],\t/a/regfile/regfile$16$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b517|t/a/regfile/reg0_b530  (
    .a({\t/a/ID_rs1 [0],_al_u803_o}),
    .b(\t/a/ID_rs1 [1:0]),
    .c({\t/a/regfile/regfile$16$ [5],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [5],\t/a/regfile/regfile$16$ [18]}),
    .e({open_n26740,\t/a/regfile/regfile$17$ [18]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u430_o,_al_u804_o}),
    .q({\t/a/regfile/regfile$16$ [5],\t/a/regfile/regfile$16$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b518|t/a/regfile/reg0_b528  (
    .a({\t/a/ID_rs1 [0],_al_u845_o}),
    .b(\t/a/ID_rs1 [1:0]),
    .c({\t/a/regfile/regfile$16$ [6],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [6],\t/a/regfile/regfile$16$ [16]}),
    .e({open_n26756,\t/a/regfile/regfile$17$ [16]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u409_o,_al_u846_o}),
    .q({\t/a/regfile/regfile$16$ [6],\t/a/regfile/regfile$16$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b519|t/a/regfile/reg0_b525  (
    .a({_al_u383_o,_al_u908_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$16$ [7],\t/a/regfile/regfile$16$ [13]}),
    .e({\t/a/regfile/regfile$17$ [7],\t/a/regfile/regfile$17$ [13]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u384_o,_al_u909_o}),
    .q({\t/a/regfile/regfile$16$ [7],\t/a/regfile/regfile$16$ [13]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b520|t/a/regfile/reg0_b523  (
    .a({\t/a/ID_rs1 [0],_al_u950_o}),
    .b(\t/a/ID_rs1 [1:0]),
    .c({\t/a/regfile/regfile$16$ [8],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [8],\t/a/regfile/regfile$16$ [11]}),
    .e({open_n26787,\t/a/regfile/regfile$17$ [11]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [11]}),
    .sr(rst_pad),
    .f({_al_u367_o,_al_u951_o}),
    .q({\t/a/regfile/regfile$16$ [8],\t/a/regfile/regfile$16$ [11]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b522|t/a/regfile/reg0_b521  (
    .a({\t/a/ID_rs1 [0],_al_u341_o}),
    .b(\t/a/ID_rs1 [1:0]),
    .c({\t/a/regfile/regfile$16$ [10],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [10],\t/a/regfile/regfile$16$ [9]}),
    .e({open_n26803,\t/a/regfile/regfile$17$ [9]}),
    .mi(\t/a/reg_writedat [10:9]),
    .sr(rst_pad),
    .f({_al_u976_o,_al_u342_o}),
    .q(\t/a/regfile/regfile$16$ [10:9]));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b524|t/a/regfile/reg0_b542  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$16$ [12],\t/a/regfile/regfile$16$ [30]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [12],\t/a/regfile/regfile$17$ [30]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u934_o,_al_u514_o}),
    .q({\t/a/regfile/regfile$16$ [12],\t/a/regfile/regfile$16$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b526|t/a/regfile/reg0_b540  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$16$ [14],\t/a/regfile/regfile$16$ [28]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [14],\t/a/regfile/regfile$17$ [28]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u892_o,_al_u577_o}),
    .q({\t/a/regfile/regfile$16$ [14],\t/a/regfile/regfile$16$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b527|t/a/regfile/reg0_b538  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$16$ [15],\t/a/regfile/regfile$16$ [26]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [15],\t/a/regfile/regfile$17$ [26]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u871_o,_al_u619_o}),
    .q({\t/a/regfile/regfile$16$ [15],\t/a/regfile/regfile$16$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b529|t/a/regfile/reg0_b537  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$16$ [17],\t/a/regfile/regfile$16$ [25]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [17],\t/a/regfile/regfile$17$ [25]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u829_o,_al_u640_o}),
    .q({\t/a/regfile/regfile$16$ [17],\t/a/regfile/regfile$16$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b531|t/a/regfile/reg0_b536  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$16$ [19],\t/a/regfile/regfile$16$ [24]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [19],\t/a/regfile/regfile$17$ [24]}),
    .mi({\t/a/reg_writedat [19],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u787_o,_al_u661_o}),
    .q({\t/a/regfile/regfile$16$ [19],\t/a/regfile/regfile$16$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b533|t/a/regfile/reg0_b535  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$16$ [21],\t/a/regfile/regfile$16$ [23]}),
    .ce(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [21],\t/a/regfile/regfile$17$ [23]}),
    .mi({\t/a/reg_writedat [21],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u724_o,_al_u682_o}),
    .q({\t/a/regfile/regfile$16$ [21],\t/a/regfile/regfile$16$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~0*~D*~C*B*A)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~1*~D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b544|t/a/regfile/reg0_b574  (
    .a({_al_u256_o,_al_u1225_o}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$16$ [30]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$17$ [30]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b544_sel_is_3_o ,_al_u1226_o}),
    .q({\t/a/regfile/regfile$17$ [0],\t/a/regfile/regfile$17$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b545|t/a/regfile/reg0_b572  (
    .a({\t/a/ID_rs2 [0],_al_u1288_o}),
    .b(\t/a/ID_rs2 [1:0]),
    .c({\t/a/regfile/regfile$16$ [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [1],\t/a/regfile/regfile$16$ [28]}),
    .e({open_n26912,\t/a/regfile/regfile$17$ [28]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1482_o,_al_u1289_o}),
    .q({\t/a/regfile/regfile$17$ [1],\t/a/regfile/regfile$17$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b546|t/a/regfile/reg0_b570  (
    .a({\t/a/ID_rs2 [0],_al_u1330_o}),
    .b(\t/a/ID_rs2 [1:0]),
    .c({\t/a/regfile/regfile$16$ [2],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [2],\t/a/regfile/regfile$16$ [26]}),
    .e({open_n26928,\t/a/regfile/regfile$17$ [26]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1251_o,_al_u1331_o}),
    .q({\t/a/regfile/regfile$17$ [2],\t/a/regfile/regfile$17$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b547|t/a/regfile/reg0_b567  (
    .a({_al_u1183_o,_al_u1393_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$16$ [3],\t/a/regfile/regfile$16$ [23]}),
    .e({\t/a/regfile/regfile$17$ [3],\t/a/regfile/regfile$17$ [23]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1184_o,_al_u1394_o}),
    .q({\t/a/regfile/regfile$17$ [3],\t/a/regfile/regfile$17$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b548|t/a/regfile/reg0_b565  (
    .a({\t/a/ID_rs2 [0],_al_u1435_o}),
    .b(\t/a/ID_rs2 [1:0]),
    .c({\t/a/regfile/regfile$16$ [4],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [4],\t/a/regfile/regfile$16$ [21]}),
    .e({open_n26959,\t/a/regfile/regfile$17$ [21]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1167_o,_al_u1436_o}),
    .q({\t/a/regfile/regfile$17$ [4],\t/a/regfile/regfile$17$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b549|t/a/regfile/reg0_b561  (
    .a({\t/a/ID_rs2 [0],_al_u1540_o}),
    .b(\t/a/ID_rs2 [1:0]),
    .c({\t/a/regfile/regfile$16$ [5],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [5],\t/a/regfile/regfile$16$ [17]}),
    .e({open_n26975,\t/a/regfile/regfile$17$ [17]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1146_o,_al_u1541_o}),
    .q({\t/a/regfile/regfile$17$ [5],\t/a/regfile/regfile$17$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b550|t/a/regfile/reg0_b559  (
    .a({\t/a/ID_rs2 [0],_al_u1582_o}),
    .b(\t/a/ID_rs2 [1:0]),
    .c({\t/a/regfile/regfile$16$ [6],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [6],\t/a/regfile/regfile$16$ [15]}),
    .e({open_n26991,\t/a/regfile/regfile$17$ [15]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u1125_o,_al_u1583_o}),
    .q({\t/a/regfile/regfile$17$ [6],\t/a/regfile/regfile$17$ [15]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b551|t/a/regfile/reg0_b556  (
    .a({\t/a/ID_rs2 [0],_al_u1645_o}),
    .b(\t/a/ID_rs2 [1:0]),
    .c({\t/a/regfile/regfile$16$ [7],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [7],\t/a/regfile/regfile$16$ [12]}),
    .e({open_n27007,\t/a/regfile/regfile$17$ [12]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u1104_o,_al_u1646_o}),
    .q({\t/a/regfile/regfile$17$ [7],\t/a/regfile/regfile$17$ [12]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b552|t/a/regfile/reg0_b554  (
    .a({_al_u1078_o,_al_u1687_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$16$ [8],\t/a/regfile/regfile$16$ [10]}),
    .e({\t/a/regfile/regfile$17$ [8],\t/a/regfile/regfile$17$ [10]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [10]}),
    .sr(rst_pad),
    .f({_al_u1079_o,_al_u1688_o}),
    .q({\t/a/regfile/regfile$17$ [8],\t/a/regfile/regfile$17$ [10]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b553|t/a/regfile/reg0_b575  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$16$ [9],\t/a/regfile/regfile$16$ [31]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [9],\t/a/regfile/regfile$17$ [31]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1062_o,_al_u1209_o}),
    .q({\t/a/regfile/regfile$17$ [9],\t/a/regfile/regfile$17$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b555|t/a/regfile/reg0_b573  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$16$ [11],\t/a/regfile/regfile$16$ [29]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [11],\t/a/regfile/regfile$17$ [29]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1671_o,_al_u1272_o}),
    .q({\t/a/regfile/regfile$17$ [11],\t/a/regfile/regfile$17$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b557|t/a/regfile/reg0_b571  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$16$ [13],\t/a/regfile/regfile$16$ [27]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [13],\t/a/regfile/regfile$17$ [27]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1629_o,_al_u1314_o}),
    .q({\t/a/regfile/regfile$17$ [13],\t/a/regfile/regfile$17$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b558|t/a/regfile/reg0_b569  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$16$ [14],\t/a/regfile/regfile$16$ [25]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [14],\t/a/regfile/regfile$17$ [25]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1608_o,_al_u1356_o}),
    .q({\t/a/regfile/regfile$17$ [14],\t/a/regfile/regfile$17$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b560|t/a/regfile/reg0_b568  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$16$ [16],\t/a/regfile/regfile$16$ [24]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [16],\t/a/regfile/regfile$17$ [24]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1566_o,_al_u1377_o}),
    .q({\t/a/regfile/regfile$17$ [16],\t/a/regfile/regfile$17$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b562|t/a/regfile/reg0_b566  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$16$ [18],\t/a/regfile/regfile$16$ [22]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [18],\t/a/regfile/regfile$17$ [22]}),
    .mi({\t/a/reg_writedat [18],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1524_o,_al_u1419_o}),
    .q({\t/a/regfile/regfile$17$ [18],\t/a/regfile/regfile$17$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b563|t/a/regfile/reg0_b564  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$16$ [19],\t/a/regfile/regfile$16$ [20]}),
    .ce(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$17$ [19],\t/a/regfile/regfile$17$ [20]}),
    .mi({\t/a/reg_writedat [19],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1503_o,_al_u1461_o}),
    .q({\t/a/regfile/regfile$17$ [19],\t/a/regfile/regfile$17$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~0*~D*C*~B*A)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~1*~D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000000100000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b576|t/a/regfile/reg0_b607  (
    .a({_al_u256_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$18$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$19$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b576_sel_is_3_o ,_al_u488_o}),
    .q({\t/a/regfile/regfile$18$ [0],\t/a/regfile/regfile$18$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b577|t/a/regfile/reg0_b592  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$18$ [1],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [1],\t/a/regfile/regfile$18$ [16]}),
    .e({open_n27144,\t/a/regfile/regfile$19$ [16]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u767_o,_al_u845_o}),
    .q({\t/a/regfile/regfile$18$ [1],\t/a/regfile/regfile$18$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b578|t/a/regfile/reg0_b606  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$18$ [2],\t/a/regfile/regfile$18$ [30]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [2],\t/a/regfile/regfile$19$ [30]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u536_o,_al_u515_o}),
    .q({\t/a/regfile/regfile$18$ [2],\t/a/regfile/regfile$18$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b579|t/a/regfile/reg0_b604  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$18$ [3],\t/a/regfile/regfile$18$ [28]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [3],\t/a/regfile/regfile$19$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u473_o,_al_u578_o}),
    .q({\t/a/regfile/regfile$18$ [3],\t/a/regfile/regfile$18$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b580|t/a/regfile/reg0_b605  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [4],\t/a/regfile/regfile$18$ [29]}),
    .e({\t/a/regfile/regfile$19$ [4],\t/a/regfile/regfile$19$ [29]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u446_o,_al_u551_o}),
    .q({\t/a/regfile/regfile$18$ [4],\t/a/regfile/regfile$18$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b581|t/a/regfile/reg0_b602  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$18$ [5],\t/a/regfile/regfile$18$ [26]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [5],\t/a/regfile/regfile$19$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u431_o,_al_u620_o}),
    .q({\t/a/regfile/regfile$18$ [5],\t/a/regfile/regfile$18$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b582|t/a/regfile/reg0_b601  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$18$ [6],\t/a/regfile/regfile$18$ [25]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [6],\t/a/regfile/regfile$19$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u410_o,_al_u641_o}),
    .q({\t/a/regfile/regfile$18$ [6],\t/a/regfile/regfile$18$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b583|t/a/regfile/reg0_b603  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [7],\t/a/regfile/regfile$18$ [27]}),
    .e({\t/a/regfile/regfile$19$ [7],\t/a/regfile/regfile$19$ [27]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u383_o,_al_u593_o}),
    .q({\t/a/regfile/regfile$18$ [7],\t/a/regfile/regfile$18$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b584|t/a/regfile/reg0_b600  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$18$ [8],\t/a/regfile/regfile$18$ [24]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [8],\t/a/regfile/regfile$19$ [24]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u368_o,_al_u662_o}),
    .q({\t/a/regfile/regfile$18$ [8],\t/a/regfile/regfile$18$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b585|t/a/regfile/reg0_b598  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [9],\t/a/regfile/regfile$18$ [22]}),
    .e({\t/a/regfile/regfile$19$ [9],\t/a/regfile/regfile$19$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u341_o,_al_u698_o}),
    .q({\t/a/regfile/regfile$18$ [9],\t/a/regfile/regfile$18$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b586|t/a/regfile/reg0_b599  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$18$ [10],\t/a/regfile/regfile$18$ [23]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [10],\t/a/regfile/regfile$19$ [23]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u977_o,_al_u683_o}),
    .q({\t/a/regfile/regfile$18$ [10],\t/a/regfile/regfile$18$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b587|t/a/regfile/reg0_b596  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [11],\t/a/regfile/regfile$18$ [20]}),
    .e({\t/a/regfile/regfile$19$ [11],\t/a/regfile/regfile$19$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u950_o,_al_u740_o}),
    .q({\t/a/regfile/regfile$18$ [11],\t/a/regfile/regfile$18$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b588|t/a/regfile/reg0_b597  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$18$ [12],\t/a/regfile/regfile$18$ [21]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [12],\t/a/regfile/regfile$19$ [21]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u935_o,_al_u725_o}),
    .q({\t/a/regfile/regfile$18$ [12],\t/a/regfile/regfile$18$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b589|t/a/regfile/reg0_b594  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [13],\t/a/regfile/regfile$18$ [18]}),
    .e({\t/a/regfile/regfile$19$ [13],\t/a/regfile/regfile$19$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u908_o,_al_u803_o}),
    .q({\t/a/regfile/regfile$18$ [13],\t/a/regfile/regfile$18$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b590|t/a/regfile/reg0_b595  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$18$ [14],\t/a/regfile/regfile$18$ [19]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [14],\t/a/regfile/regfile$19$ [19]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u893_o,_al_u788_o}),
    .q({\t/a/regfile/regfile$18$ [14],\t/a/regfile/regfile$18$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b591|t/a/regfile/reg0_b593  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$18$ [15],\t/a/regfile/regfile$18$ [17]}),
    .ce(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [15],\t/a/regfile/regfile$19$ [17]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u872_o,_al_u830_o}),
    .q({\t/a/regfile/regfile$18$ [15],\t/a/regfile/regfile$18$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~0*~D*C*B*A)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~1*~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b608|t/a/regfile/reg0_b638  (
    .a({_al_u256_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$18$ [30]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$19$ [30]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b608_sel_is_3_o ,_al_u1225_o}),
    .q({\t/a/regfile/regfile$19$ [0],\t/a/regfile/regfile$19$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b609|t/a/regfile/reg0_b639  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$18$ [1],\t/a/regfile/regfile$18$ [31]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [1],\t/a/regfile/regfile$19$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1483_o,_al_u1210_o}),
    .q({\t/a/regfile/regfile$19$ [1],\t/a/regfile/regfile$19$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b610|t/a/regfile/reg0_b637  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$18$ [2],\t/a/regfile/regfile$18$ [29]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [2],\t/a/regfile/regfile$19$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1252_o,_al_u1273_o}),
    .q({\t/a/regfile/regfile$19$ [2],\t/a/regfile/regfile$19$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b611|t/a/regfile/reg0_b636  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [3],\t/a/regfile/regfile$18$ [28]}),
    .e({\t/a/regfile/regfile$19$ [3],\t/a/regfile/regfile$19$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1183_o,_al_u1288_o}),
    .q({\t/a/regfile/regfile$19$ [3],\t/a/regfile/regfile$19$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b612|t/a/regfile/reg0_b635  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$18$ [4],\t/a/regfile/regfile$18$ [27]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [4],\t/a/regfile/regfile$19$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1168_o,_al_u1315_o}),
    .q({\t/a/regfile/regfile$19$ [4],\t/a/regfile/regfile$19$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b613|t/a/regfile/reg0_b633  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$18$ [5],\t/a/regfile/regfile$18$ [25]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [5],\t/a/regfile/regfile$19$ [25]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1147_o,_al_u1357_o}),
    .q({\t/a/regfile/regfile$19$ [5],\t/a/regfile/regfile$19$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b614|t/a/regfile/reg0_b632  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$18$ [6],\t/a/regfile/regfile$18$ [24]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [6],\t/a/regfile/regfile$19$ [24]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1126_o,_al_u1378_o}),
    .q({\t/a/regfile/regfile$19$ [6],\t/a/regfile/regfile$19$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b615|t/a/regfile/reg0_b630  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$18$ [7],\t/a/regfile/regfile$18$ [22]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [7],\t/a/regfile/regfile$19$ [22]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1105_o,_al_u1420_o}),
    .q({\t/a/regfile/regfile$19$ [7],\t/a/regfile/regfile$19$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b616|t/a/regfile/reg0_b634  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [8],\t/a/regfile/regfile$18$ [26]}),
    .e({\t/a/regfile/regfile$19$ [8],\t/a/regfile/regfile$19$ [26]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1078_o,_al_u1330_o}),
    .q({\t/a/regfile/regfile$19$ [8],\t/a/regfile/regfile$19$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b617|t/a/regfile/reg0_b628  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$18$ [9],\t/a/regfile/regfile$18$ [20]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [9],\t/a/regfile/regfile$19$ [20]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1063_o,_al_u1462_o}),
    .q({\t/a/regfile/regfile$19$ [9],\t/a/regfile/regfile$19$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b618|t/a/regfile/reg0_b631  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [10],\t/a/regfile/regfile$18$ [23]}),
    .e({\t/a/regfile/regfile$19$ [10],\t/a/regfile/regfile$19$ [23]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1687_o,_al_u1393_o}),
    .q({\t/a/regfile/regfile$19$ [10],\t/a/regfile/regfile$19$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b619|t/a/regfile/reg0_b627  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$18$ [11],\t/a/regfile/regfile$18$ [19]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [11],\t/a/regfile/regfile$19$ [19]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1672_o,_al_u1504_o}),
    .q({\t/a/regfile/regfile$19$ [11],\t/a/regfile/regfile$19$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b620|t/a/regfile/reg0_b629  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [12],\t/a/regfile/regfile$18$ [21]}),
    .e({\t/a/regfile/regfile$19$ [12],\t/a/regfile/regfile$19$ [21]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1645_o,_al_u1435_o}),
    .q({\t/a/regfile/regfile$19$ [12],\t/a/regfile/regfile$19$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b621|t/a/regfile/reg0_b626  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$18$ [13],\t/a/regfile/regfile$18$ [18]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [13],\t/a/regfile/regfile$19$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1630_o,_al_u1525_o}),
    .q({\t/a/regfile/regfile$19$ [13],\t/a/regfile/regfile$19$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b622|t/a/regfile/reg0_b624  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$18$ [14],\t/a/regfile/regfile$18$ [16]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$19$ [14],\t/a/regfile/regfile$19$ [16]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1609_o,_al_u1567_o}),
    .q({\t/a/regfile/regfile$19$ [14],\t/a/regfile/regfile$19$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b623|t/a/regfile/reg0_b625  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$18$ [15],\t/a/regfile/regfile$18$ [17]}),
    .e({\t/a/regfile/regfile$19$ [15],\t/a/regfile/regfile$19$ [17]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1582_o,_al_u1540_o}),
    .q({\t/a/regfile/regfile$19$ [15],\t/a/regfile/regfile$19$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b641|t/a/regfile/reg0_b670  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$20$ [1],\t/a/regfile/regfile$20$ [30]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [1],\t/a/regfile/regfile$21$ [30]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u764_o,_al_u512_o}),
    .q({\t/a/regfile/regfile$20$ [1],\t/a/regfile/regfile$20$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b642|t/a/regfile/reg0_b668  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$20$ [2],\t/a/regfile/regfile$20$ [28]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [2],\t/a/regfile/regfile$21$ [28]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u533_o,_al_u575_o}),
    .q({\t/a/regfile/regfile$20$ [2],\t/a/regfile/regfile$20$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b643|t/a/regfile/reg0_b666  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$20$ [3],\t/a/regfile/regfile$20$ [26]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [3],\t/a/regfile/regfile$21$ [26]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u470_o,_al_u617_o}),
    .q({\t/a/regfile/regfile$20$ [3],\t/a/regfile/regfile$20$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b645|t/a/regfile/reg0_b665  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$20$ [5],\t/a/regfile/regfile$20$ [25]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [5],\t/a/regfile/regfile$21$ [25]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u428_o,_al_u638_o}),
    .q({\t/a/regfile/regfile$20$ [5],\t/a/regfile/regfile$20$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b646|t/a/regfile/reg0_b664  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$20$ [6],\t/a/regfile/regfile$20$ [24]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [6],\t/a/regfile/regfile$21$ [24]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u407_o,_al_u659_o}),
    .q({\t/a/regfile/regfile$20$ [6],\t/a/regfile/regfile$20$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b648|t/a/regfile/reg0_b663  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$20$ [8],\t/a/regfile/regfile$20$ [23]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [8],\t/a/regfile/regfile$21$ [23]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u365_o,_al_u680_o}),
    .q({\t/a/regfile/regfile$20$ [8],\t/a/regfile/regfile$20$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b650|t/a/regfile/reg0_b661  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$20$ [10],\t/a/regfile/regfile$20$ [21]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [10],\t/a/regfile/regfile$21$ [21]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u974_o,_al_u722_o}),
    .q({\t/a/regfile/regfile$20$ [10],\t/a/regfile/regfile$20$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b652|t/a/regfile/reg0_b659  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$20$ [12],\t/a/regfile/regfile$20$ [19]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [12],\t/a/regfile/regfile$21$ [19]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u932_o,_al_u785_o}),
    .q({\t/a/regfile/regfile$20$ [12],\t/a/regfile/regfile$20$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b654|t/a/regfile/reg0_b657  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$20$ [14],\t/a/regfile/regfile$20$ [17]}),
    .ce(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [14],\t/a/regfile/regfile$21$ [17]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u890_o,_al_u827_o}),
    .q({\t/a/regfile/regfile$20$ [14],\t/a/regfile/regfile$20$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b65|t/a/regfile/reg0_b68  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$2$ [1],\t/a/regfile/regfile$3$ [4]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$3$ [1],\t/a/regfile/regfile$2$ [4]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [4]}),
    .sr(rst_pad),
    .f({_al_u757_o,_al_u452_o}),
    .q({\t/a/regfile/regfile$2$ [1],\t/a/regfile/regfile$2$ [4]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b66|t/a/regfile/reg0_b67  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$2$ [2],\t/a/regfile/regfile$2$ [3]}),
    .ce(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$3$ [2],\t/a/regfile/regfile$3$ [3]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u526_o,_al_u463_o}),
    .q({\t/a/regfile/regfile$2$ [2],\t/a/regfile/regfile$2$ [3]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b673|t/a/regfile/reg0_b703  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$20$ [1],\t/a/regfile/regfile$20$ [31]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [1],\t/a/regfile/regfile$21$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1480_o,_al_u1207_o}),
    .q({\t/a/regfile/regfile$21$ [1],\t/a/regfile/regfile$21$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b674|t/a/regfile/reg0_b701  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$20$ [2],\t/a/regfile/regfile$20$ [29]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [2],\t/a/regfile/regfile$21$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1249_o,_al_u1270_o}),
    .q({\t/a/regfile/regfile$21$ [2],\t/a/regfile/regfile$21$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b676|t/a/regfile/reg0_b699  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$20$ [4],\t/a/regfile/regfile$20$ [27]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [4],\t/a/regfile/regfile$21$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1165_o,_al_u1312_o}),
    .q({\t/a/regfile/regfile$21$ [4],\t/a/regfile/regfile$21$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b677|t/a/regfile/reg0_b697  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$20$ [5],\t/a/regfile/regfile$20$ [25]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [5],\t/a/regfile/regfile$21$ [25]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1144_o,_al_u1354_o}),
    .q({\t/a/regfile/regfile$21$ [5],\t/a/regfile/regfile$21$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b678|t/a/regfile/reg0_b696  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$20$ [6],\t/a/regfile/regfile$20$ [24]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [6],\t/a/regfile/regfile$21$ [24]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1123_o,_al_u1375_o}),
    .q({\t/a/regfile/regfile$21$ [6],\t/a/regfile/regfile$21$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b679|t/a/regfile/reg0_b694  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$20$ [7],\t/a/regfile/regfile$20$ [22]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [7],\t/a/regfile/regfile$21$ [22]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1102_o,_al_u1417_o}),
    .q({\t/a/regfile/regfile$21$ [7],\t/a/regfile/regfile$21$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b681|t/a/regfile/reg0_b692  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$20$ [9],\t/a/regfile/regfile$20$ [20]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [9],\t/a/regfile/regfile$21$ [20]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1060_o,_al_u1459_o}),
    .q({\t/a/regfile/regfile$21$ [9],\t/a/regfile/regfile$21$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b683|t/a/regfile/reg0_b691  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$20$ [11],\t/a/regfile/regfile$20$ [19]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [11],\t/a/regfile/regfile$21$ [19]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1669_o,_al_u1501_o}),
    .q({\t/a/regfile/regfile$21$ [11],\t/a/regfile/regfile$21$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b685|t/a/regfile/reg0_b690  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$20$ [13],\t/a/regfile/regfile$20$ [18]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [13],\t/a/regfile/regfile$21$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1627_o,_al_u1522_o}),
    .q({\t/a/regfile/regfile$21$ [13],\t/a/regfile/regfile$21$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b686|t/a/regfile/reg0_b688  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$20$ [14],\t/a/regfile/regfile$20$ [16]}),
    .ce(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$21$ [14],\t/a/regfile/regfile$21$ [16]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1606_o,_al_u1564_o}),
    .q({\t/a/regfile/regfile$21$ [14],\t/a/regfile/regfile$21$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~0*D*C*~B*A)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~1*D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b704|t/a/regfile/reg0_b735  (
    .a({_al_u256_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$22$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$23$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b704_sel_is_3_o ,_al_u486_o}),
    .q({\t/a/regfile/regfile$22$ [0],\t/a/regfile/regfile$22$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b705|t/a/regfile/reg0_b720  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$22$ [1],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [1],\t/a/regfile/regfile$22$ [16]}),
    .e({open_n27860,\t/a/regfile/regfile$23$ [16]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u765_o,_al_u843_o}),
    .q({\t/a/regfile/regfile$22$ [1],\t/a/regfile/regfile$22$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b706|t/a/regfile/reg0_b734  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$22$ [2],\t/a/regfile/regfile$22$ [30]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [2],\t/a/regfile/regfile$23$ [30]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u534_o,_al_u513_o}),
    .q({\t/a/regfile/regfile$22$ [2],\t/a/regfile/regfile$22$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b707|t/a/regfile/reg0_b732  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$22$ [3],\t/a/regfile/regfile$22$ [28]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [3],\t/a/regfile/regfile$23$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u471_o,_al_u576_o}),
    .q({\t/a/regfile/regfile$22$ [3],\t/a/regfile/regfile$22$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b708|t/a/regfile/reg0_b733  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [4],\t/a/regfile/regfile$22$ [29]}),
    .e({\t/a/regfile/regfile$23$ [4],\t/a/regfile/regfile$23$ [29]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u444_o,_al_u549_o}),
    .q({\t/a/regfile/regfile$22$ [4],\t/a/regfile/regfile$22$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b709|t/a/regfile/reg0_b730  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$22$ [5],\t/a/regfile/regfile$22$ [26]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [5],\t/a/regfile/regfile$23$ [26]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u429_o,_al_u618_o}),
    .q({\t/a/regfile/regfile$22$ [5],\t/a/regfile/regfile$22$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b710|t/a/regfile/reg0_b729  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$22$ [6],\t/a/regfile/regfile$22$ [25]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [6],\t/a/regfile/regfile$23$ [25]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u408_o,_al_u639_o}),
    .q({\t/a/regfile/regfile$22$ [6],\t/a/regfile/regfile$22$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b711|t/a/regfile/reg0_b731  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [7],\t/a/regfile/regfile$22$ [27]}),
    .e({\t/a/regfile/regfile$23$ [7],\t/a/regfile/regfile$23$ [27]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u381_o,_al_u591_o}),
    .q({\t/a/regfile/regfile$22$ [7],\t/a/regfile/regfile$22$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b712|t/a/regfile/reg0_b728  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$22$ [8],\t/a/regfile/regfile$22$ [24]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [8],\t/a/regfile/regfile$23$ [24]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u366_o,_al_u660_o}),
    .q({\t/a/regfile/regfile$22$ [8],\t/a/regfile/regfile$22$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b713|t/a/regfile/reg0_b726  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [9],\t/a/regfile/regfile$22$ [22]}),
    .e({\t/a/regfile/regfile$23$ [9],\t/a/regfile/regfile$23$ [22]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u339_o,_al_u696_o}),
    .q({\t/a/regfile/regfile$22$ [9],\t/a/regfile/regfile$22$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b714|t/a/regfile/reg0_b727  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$22$ [10],\t/a/regfile/regfile$22$ [23]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [10],\t/a/regfile/regfile$23$ [23]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u975_o,_al_u681_o}),
    .q({\t/a/regfile/regfile$22$ [10],\t/a/regfile/regfile$22$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b715|t/a/regfile/reg0_b724  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [11],\t/a/regfile/regfile$22$ [20]}),
    .e({\t/a/regfile/regfile$23$ [11],\t/a/regfile/regfile$23$ [20]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u948_o,_al_u738_o}),
    .q({\t/a/regfile/regfile$22$ [11],\t/a/regfile/regfile$22$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b716|t/a/regfile/reg0_b725  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$22$ [12],\t/a/regfile/regfile$22$ [21]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [12],\t/a/regfile/regfile$23$ [21]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u933_o,_al_u723_o}),
    .q({\t/a/regfile/regfile$22$ [12],\t/a/regfile/regfile$22$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b717|t/a/regfile/reg0_b722  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [13],\t/a/regfile/regfile$22$ [18]}),
    .e({\t/a/regfile/regfile$23$ [13],\t/a/regfile/regfile$23$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u906_o,_al_u801_o}),
    .q({\t/a/regfile/regfile$22$ [13],\t/a/regfile/regfile$22$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b718|t/a/regfile/reg0_b723  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$22$ [14],\t/a/regfile/regfile$22$ [19]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [14],\t/a/regfile/regfile$23$ [19]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u891_o,_al_u786_o}),
    .q({\t/a/regfile/regfile$22$ [14],\t/a/regfile/regfile$22$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b719|t/a/regfile/reg0_b721  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$22$ [15],\t/a/regfile/regfile$22$ [17]}),
    .ce(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [15],\t/a/regfile/regfile$23$ [17]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u870_o,_al_u828_o}),
    .q({\t/a/regfile/regfile$22$ [15],\t/a/regfile/regfile$22$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~0*D*C*B*A)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~1*D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b736|t/a/regfile/reg0_b766  (
    .a({_al_u256_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$22$ [30]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$23$ [30]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b736_sel_is_3_o ,_al_u1223_o}),
    .q({\t/a/regfile/regfile$23$ [0],\t/a/regfile/regfile$23$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b737|t/a/regfile/reg0_b767  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$22$ [1],\t/a/regfile/regfile$22$ [31]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [1],\t/a/regfile/regfile$23$ [31]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u1481_o,_al_u1208_o}),
    .q({\t/a/regfile/regfile$23$ [1],\t/a/regfile/regfile$23$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b738|t/a/regfile/reg0_b765  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$22$ [2],\t/a/regfile/regfile$22$ [29]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [2],\t/a/regfile/regfile$23$ [29]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1250_o,_al_u1271_o}),
    .q({\t/a/regfile/regfile$23$ [2],\t/a/regfile/regfile$23$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b739|t/a/regfile/reg0_b764  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [3],\t/a/regfile/regfile$22$ [28]}),
    .e({\t/a/regfile/regfile$23$ [3],\t/a/regfile/regfile$23$ [28]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1181_o,_al_u1286_o}),
    .q({\t/a/regfile/regfile$23$ [3],\t/a/regfile/regfile$23$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b740|t/a/regfile/reg0_b763  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$22$ [4],\t/a/regfile/regfile$22$ [27]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [4],\t/a/regfile/regfile$23$ [27]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1166_o,_al_u1313_o}),
    .q({\t/a/regfile/regfile$23$ [4],\t/a/regfile/regfile$23$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b741|t/a/regfile/reg0_b761  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$22$ [5],\t/a/regfile/regfile$22$ [25]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [5],\t/a/regfile/regfile$23$ [25]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1145_o,_al_u1355_o}),
    .q({\t/a/regfile/regfile$23$ [5],\t/a/regfile/regfile$23$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b742|t/a/regfile/reg0_b760  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$22$ [6],\t/a/regfile/regfile$22$ [24]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [6],\t/a/regfile/regfile$23$ [24]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1124_o,_al_u1376_o}),
    .q({\t/a/regfile/regfile$23$ [6],\t/a/regfile/regfile$23$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b743|t/a/regfile/reg0_b758  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$22$ [7],\t/a/regfile/regfile$22$ [22]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [7],\t/a/regfile/regfile$23$ [22]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1103_o,_al_u1418_o}),
    .q({\t/a/regfile/regfile$23$ [7],\t/a/regfile/regfile$23$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b744|t/a/regfile/reg0_b762  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [8],\t/a/regfile/regfile$22$ [26]}),
    .e({\t/a/regfile/regfile$23$ [8],\t/a/regfile/regfile$23$ [26]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1076_o,_al_u1328_o}),
    .q({\t/a/regfile/regfile$23$ [8],\t/a/regfile/regfile$23$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b745|t/a/regfile/reg0_b756  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$22$ [9],\t/a/regfile/regfile$22$ [20]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [9],\t/a/regfile/regfile$23$ [20]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1061_o,_al_u1460_o}),
    .q({\t/a/regfile/regfile$23$ [9],\t/a/regfile/regfile$23$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b746|t/a/regfile/reg0_b759  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [10],\t/a/regfile/regfile$22$ [23]}),
    .e({\t/a/regfile/regfile$23$ [10],\t/a/regfile/regfile$23$ [23]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1685_o,_al_u1391_o}),
    .q({\t/a/regfile/regfile$23$ [10],\t/a/regfile/regfile$23$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b747|t/a/regfile/reg0_b755  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$22$ [11],\t/a/regfile/regfile$22$ [19]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [11],\t/a/regfile/regfile$23$ [19]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1670_o,_al_u1502_o}),
    .q({\t/a/regfile/regfile$23$ [11],\t/a/regfile/regfile$23$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b748|t/a/regfile/reg0_b757  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [12],\t/a/regfile/regfile$22$ [21]}),
    .e({\t/a/regfile/regfile$23$ [12],\t/a/regfile/regfile$23$ [21]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1643_o,_al_u1433_o}),
    .q({\t/a/regfile/regfile$23$ [12],\t/a/regfile/regfile$23$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b749|t/a/regfile/reg0_b754  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$22$ [13],\t/a/regfile/regfile$22$ [18]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [13],\t/a/regfile/regfile$23$ [18]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1628_o,_al_u1523_o}),
    .q({\t/a/regfile/regfile$23$ [13],\t/a/regfile/regfile$23$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b750|t/a/regfile/reg0_b752  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$22$ [14],\t/a/regfile/regfile$22$ [16]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$23$ [14],\t/a/regfile/regfile$23$ [16]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1607_o,_al_u1565_o}),
    .q({\t/a/regfile/regfile$23$ [14],\t/a/regfile/regfile$23$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b751|t/a/regfile/reg0_b753  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$22$ [15],\t/a/regfile/regfile$22$ [17]}),
    .e({\t/a/regfile/regfile$23$ [15],\t/a/regfile/regfile$23$ [17]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u1580_o,_al_u1538_o}),
    .q({\t/a/regfile/regfile$23$ [15],\t/a/regfile/regfile$23$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b768|t/a/regfile/reg0_b798  (
    .a({_al_u256_o,_al_u519_o}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$24$ [30]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$25$ [30]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b768_sel_is_3_o ,_al_u520_o}),
    .q({\t/a/regfile/regfile$24$ [0],\t/a/regfile/regfile$24$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b769|t/a/regfile/reg0_b796  (
    .a({_al_u771_o,_al_u582_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [1],\t/a/regfile/regfile$24$ [28]}),
    .e({\t/a/regfile/regfile$25$ [1],\t/a/regfile/regfile$25$ [28]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u772_o,_al_u583_o}),
    .q({\t/a/regfile/regfile$24$ [1],\t/a/regfile/regfile$24$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b770|t/a/regfile/reg0_b794  (
    .a({_al_u540_o,_al_u624_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [2],\t/a/regfile/regfile$24$ [26]}),
    .e({\t/a/regfile/regfile$25$ [2],\t/a/regfile/regfile$25$ [26]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u541_o,_al_u625_o}),
    .q({\t/a/regfile/regfile$24$ [2],\t/a/regfile/regfile$24$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b771|t/a/regfile/reg0_b793  (
    .a({_al_u477_o,_al_u645_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [3],\t/a/regfile/regfile$24$ [25]}),
    .e({\t/a/regfile/regfile$25$ [3],\t/a/regfile/regfile$25$ [25]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u478_o,_al_u646_o}),
    .q({\t/a/regfile/regfile$24$ [3],\t/a/regfile/regfile$24$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b772|t/a/regfile/reg0_b792  (
    .a({\t/a/ID_rs1 [0],_al_u666_o}),
    .b(\t/a/ID_rs1 [1:0]),
    .c({\t/a/regfile/regfile$24$ [4],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [4],\t/a/regfile/regfile$24$ [24]}),
    .e({open_n28348,\t/a/regfile/regfile$25$ [24]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u441_o,_al_u667_o}),
    .q({\t/a/regfile/regfile$24$ [4],\t/a/regfile/regfile$24$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b773|t/a/regfile/reg0_b791  (
    .a({_al_u435_o,_al_u687_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [5],\t/a/regfile/regfile$24$ [23]}),
    .e({\t/a/regfile/regfile$25$ [5],\t/a/regfile/regfile$25$ [23]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u436_o,_al_u688_o}),
    .q({\t/a/regfile/regfile$24$ [5],\t/a/regfile/regfile$24$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b774|t/a/regfile/reg0_b789  (
    .a({_al_u414_o,_al_u729_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [6],\t/a/regfile/regfile$24$ [21]}),
    .e({\t/a/regfile/regfile$25$ [6],\t/a/regfile/regfile$25$ [21]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u415_o,_al_u730_o}),
    .q({\t/a/regfile/regfile$24$ [6],\t/a/regfile/regfile$24$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b775|t/a/regfile/reg0_b787  (
    .a({\t/a/ID_rs1 [0],_al_u792_o}),
    .b(\t/a/ID_rs1 [1:0]),
    .c({\t/a/regfile/regfile$24$ [7],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [7],\t/a/regfile/regfile$24$ [19]}),
    .e({open_n28394,\t/a/regfile/regfile$25$ [19]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u378_o,_al_u793_o}),
    .q({\t/a/regfile/regfile$24$ [7],\t/a/regfile/regfile$24$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b776|t/a/regfile/reg0_b785  (
    .a({_al_u372_o,_al_u834_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [8],\t/a/regfile/regfile$24$ [17]}),
    .e({\t/a/regfile/regfile$25$ [8],\t/a/regfile/regfile$25$ [17]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u373_o,_al_u835_o}),
    .q({\t/a/regfile/regfile$24$ [8],\t/a/regfile/regfile$24$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b777|t/a/regfile/reg0_b783  (
    .a({\t/a/ID_rs1 [0],_al_u876_o}),
    .b(\t/a/ID_rs1 [1:0]),
    .c({\t/a/regfile/regfile$24$ [9],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [9],\t/a/regfile/regfile$24$ [15]}),
    .e({open_n28425,\t/a/regfile/regfile$25$ [15]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u336_o,_al_u877_o}),
    .q({\t/a/regfile/regfile$24$ [9],\t/a/regfile/regfile$24$ [15]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b778|t/a/regfile/reg0_b782  (
    .a({_al_u981_o,_al_u897_o}),
    .b({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .c({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [10],\t/a/regfile/regfile$24$ [14]}),
    .e({\t/a/regfile/regfile$25$ [10],\t/a/regfile/regfile$25$ [14]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u982_o,_al_u898_o}),
    .q({\t/a/regfile/regfile$24$ [10],\t/a/regfile/regfile$24$ [14]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b779|t/a/regfile/reg0_b780  (
    .a({\t/a/ID_rs1 [0],_al_u939_o}),
    .b(\t/a/ID_rs1 [1:0]),
    .c({\t/a/regfile/regfile$24$ [11],\t/a/ID_rs1 [1]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [11],\t/a/regfile/regfile$24$ [12]}),
    .e({open_n28456,\t/a/regfile/regfile$25$ [12]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [12]}),
    .sr(rst_pad),
    .f({_al_u945_o,_al_u940_o}),
    .q({\t/a/regfile/regfile$24$ [11],\t/a/regfile/regfile$24$ [12]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b781|t/a/regfile/reg0_b799  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$24$ [13],\t/a/regfile/regfile$24$ [31]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [13],\t/a/regfile/regfile$25$ [31]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u903_o,_al_u483_o}),
    .q({\t/a/regfile/regfile$24$ [13],\t/a/regfile/regfile$24$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b784|t/a/regfile/reg0_b797  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$24$ [16],\t/a/regfile/regfile$24$ [29]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [16],\t/a/regfile/regfile$25$ [29]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u840_o,_al_u546_o}),
    .q({\t/a/regfile/regfile$24$ [16],\t/a/regfile/regfile$24$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b786|t/a/regfile/reg0_b795  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$24$ [18],\t/a/regfile/regfile$24$ [27]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [18],\t/a/regfile/regfile$25$ [27]}),
    .mi({\t/a/reg_writedat [18],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u798_o,_al_u588_o}),
    .q({\t/a/regfile/regfile$24$ [18],\t/a/regfile/regfile$24$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b788|t/a/regfile/reg0_b790  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$24$ [20],\t/a/regfile/regfile$24$ [22]}),
    .ce(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [20],\t/a/regfile/regfile$25$ [22]}),
    .mi({\t/a/reg_writedat [20],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u735_o,_al_u693_o}),
    .q({\t/a/regfile/regfile$24$ [20],\t/a/regfile/regfile$24$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(0*~D*~C*B*A)"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(1*~D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b800|t/a/regfile/reg0_b831  (
    .a({_al_u256_o,_al_u1214_o}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$24$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$25$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b800_sel_is_3_o ,_al_u1215_o}),
    .q({\t/a/regfile/regfile$25$ [0],\t/a/regfile/regfile$25$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b801|t/a/regfile/reg0_b829  (
    .a({_al_u1487_o,_al_u1277_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [1],\t/a/regfile/regfile$24$ [29]}),
    .e({\t/a/regfile/regfile$25$ [1],\t/a/regfile/regfile$25$ [29]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1488_o,_al_u1278_o}),
    .q({\t/a/regfile/regfile$25$ [1],\t/a/regfile/regfile$25$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b802|t/a/regfile/reg0_b827  (
    .a({_al_u1256_o,_al_u1319_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [2],\t/a/regfile/regfile$24$ [27]}),
    .e({\t/a/regfile/regfile$25$ [2],\t/a/regfile/regfile$25$ [27]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1257_o,_al_u1320_o}),
    .q({\t/a/regfile/regfile$25$ [2],\t/a/regfile/regfile$25$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b803|t/a/regfile/reg0_b825  (
    .a({\t/a/ID_rs2 [0],_al_u1361_o}),
    .b(\t/a/ID_rs2 [1:0]),
    .c({\t/a/regfile/regfile$24$ [3],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [3],\t/a/regfile/regfile$24$ [25]}),
    .e({open_n28569,\t/a/regfile/regfile$25$ [25]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1178_o,_al_u1362_o}),
    .q({\t/a/regfile/regfile$25$ [3],\t/a/regfile/regfile$25$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b804|t/a/regfile/reg0_b824  (
    .a({_al_u1172_o,_al_u1382_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [4],\t/a/regfile/regfile$24$ [24]}),
    .e({\t/a/regfile/regfile$25$ [4],\t/a/regfile/regfile$25$ [24]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1173_o,_al_u1383_o}),
    .q({\t/a/regfile/regfile$25$ [4],\t/a/regfile/regfile$25$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b805|t/a/regfile/reg0_b822  (
    .a({_al_u1151_o,_al_u1424_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [5],\t/a/regfile/regfile$24$ [22]}),
    .e({\t/a/regfile/regfile$25$ [5],\t/a/regfile/regfile$25$ [22]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1152_o,_al_u1425_o}),
    .q({\t/a/regfile/regfile$25$ [5],\t/a/regfile/regfile$25$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b806|t/a/regfile/reg0_b820  (
    .a({_al_u1130_o,_al_u1466_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [6],\t/a/regfile/regfile$24$ [20]}),
    .e({\t/a/regfile/regfile$25$ [6],\t/a/regfile/regfile$25$ [20]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1131_o,_al_u1467_o}),
    .q({\t/a/regfile/regfile$25$ [6],\t/a/regfile/regfile$25$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b807|t/a/regfile/reg0_b819  (
    .a({_al_u1109_o,_al_u1508_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [7],\t/a/regfile/regfile$24$ [19]}),
    .e({\t/a/regfile/regfile$25$ [7],\t/a/regfile/regfile$25$ [19]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1110_o,_al_u1509_o}),
    .q({\t/a/regfile/regfile$25$ [7],\t/a/regfile/regfile$25$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b808|t/a/regfile/reg0_b818  (
    .a({\t/a/ID_rs2 [0],_al_u1529_o}),
    .b(\t/a/ID_rs2 [1:0]),
    .c({\t/a/regfile/regfile$24$ [8],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [8],\t/a/regfile/regfile$24$ [18]}),
    .e({open_n28645,\t/a/regfile/regfile$25$ [18]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1073_o,_al_u1530_o}),
    .q({\t/a/regfile/regfile$25$ [8],\t/a/regfile/regfile$25$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b809|t/a/regfile/reg0_b816  (
    .a({_al_u1067_o,_al_u1571_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [9],\t/a/regfile/regfile$24$ [16]}),
    .e({\t/a/regfile/regfile$25$ [9],\t/a/regfile/regfile$25$ [16]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1068_o,_al_u1572_o}),
    .q({\t/a/regfile/regfile$25$ [9],\t/a/regfile/regfile$25$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b0000000100100011),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b0000000100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b810|t/a/regfile/reg0_b814  (
    .a({\t/a/ID_rs2 [0],_al_u1613_o}),
    .b(\t/a/ID_rs2 [1:0]),
    .c({\t/a/regfile/regfile$24$ [10],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [10],\t/a/regfile/regfile$24$ [14]}),
    .e({open_n28676,\t/a/regfile/regfile$25$ [14]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1682_o,_al_u1614_o}),
    .q({\t/a/regfile/regfile$25$ [10],\t/a/regfile/regfile$25$ [14]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTF1("(A*~(~C*~(D*~(0)*~(B)+D*0*~(B)+~(D)*0*B+D*0*B)))"),
    //.LUTG0("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    //.LUTG1("(A*~(~C*~(D*~(1)*~(B)+D*1*~(B)+~(D)*1*B+D*1*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010001010100000),
    .INIT_LUTF1(16'b1010001010100000),
    .INIT_LUTG0(16'b1010101010101000),
    .INIT_LUTG1(16'b1010101010101000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b811|t/a/regfile/reg0_b813  (
    .a({_al_u1676_o,_al_u1634_o}),
    .b({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .c({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$24$ [11],\t/a/regfile/regfile$24$ [13]}),
    .e({\t/a/regfile/regfile$25$ [11],\t/a/regfile/regfile$25$ [13]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [13]}),
    .sr(rst_pad),
    .f({_al_u1677_o,_al_u1635_o}),
    .q({\t/a/regfile/regfile$25$ [11],\t/a/regfile/regfile$25$ [13]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b812|t/a/regfile/reg0_b830  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$24$ [12],\t/a/regfile/regfile$24$ [30]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [12],\t/a/regfile/regfile$25$ [30]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1640_o,_al_u1220_o}),
    .q({\t/a/regfile/regfile$25$ [12],\t/a/regfile/regfile$25$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b815|t/a/regfile/reg0_b828  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$24$ [15],\t/a/regfile/regfile$24$ [28]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [15],\t/a/regfile/regfile$25$ [28]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1577_o,_al_u1283_o}),
    .q({\t/a/regfile/regfile$25$ [15],\t/a/regfile/regfile$25$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b817|t/a/regfile/reg0_b826  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$24$ [17],\t/a/regfile/regfile$24$ [26]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [17],\t/a/regfile/regfile$25$ [26]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1535_o,_al_u1325_o}),
    .q({\t/a/regfile/regfile$25$ [17],\t/a/regfile/regfile$25$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b821|t/a/regfile/reg0_b823  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$24$ [21],\t/a/regfile/regfile$24$ [23]}),
    .ce(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$25$ [21],\t/a/regfile/regfile$25$ [23]}),
    .mi({\t/a/reg_writedat [21],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1430_o,_al_u1388_o}),
    .q({\t/a/regfile/regfile$25$ [21],\t/a/regfile/regfile$25$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*~D*C*~B*A)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*~D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b832|t/a/regfile/reg0_b862  (
    .a({_al_u256_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$26$ [30]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$27$ [30]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b832_sel_is_3_o ,_al_u519_o}),
    .q({\t/a/regfile/regfile$26$ [0],\t/a/regfile/regfile$26$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b833|t/a/regfile/reg0_b860  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [1],\t/a/regfile/regfile$26$ [28]}),
    .e({\t/a/regfile/regfile$27$ [1],\t/a/regfile/regfile$27$ [28]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u771_o,_al_u582_o}),
    .q({\t/a/regfile/regfile$26$ [1],\t/a/regfile/regfile$26$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b834|t/a/regfile/reg0_b858  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [2],\t/a/regfile/regfile$26$ [26]}),
    .e({\t/a/regfile/regfile$27$ [2],\t/a/regfile/regfile$27$ [26]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u540_o,_al_u624_o}),
    .q({\t/a/regfile/regfile$26$ [2],\t/a/regfile/regfile$26$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b835|t/a/regfile/reg0_b857  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [3],\t/a/regfile/regfile$26$ [25]}),
    .e({\t/a/regfile/regfile$27$ [3],\t/a/regfile/regfile$27$ [25]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u477_o,_al_u645_o}),
    .q({\t/a/regfile/regfile$26$ [3],\t/a/regfile/regfile$26$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b836|t/a/regfile/reg0_b863  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$26$ [4],\t/a/regfile/regfile$26$ [31]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [4],\t/a/regfile/regfile$27$ [31]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u442_o,_al_u484_o}),
    .q({\t/a/regfile/regfile$26$ [4],\t/a/regfile/regfile$26$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b837|t/a/regfile/reg0_b856  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [5],\t/a/regfile/regfile$26$ [24]}),
    .e({\t/a/regfile/regfile$27$ [5],\t/a/regfile/regfile$27$ [24]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u435_o,_al_u666_o}),
    .q({\t/a/regfile/regfile$26$ [5],\t/a/regfile/regfile$26$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b838|t/a/regfile/reg0_b855  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [6],\t/a/regfile/regfile$26$ [23]}),
    .e({\t/a/regfile/regfile$27$ [6],\t/a/regfile/regfile$27$ [23]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u414_o,_al_u687_o}),
    .q({\t/a/regfile/regfile$26$ [6],\t/a/regfile/regfile$26$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b839|t/a/regfile/reg0_b861  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$26$ [7],\t/a/regfile/regfile$26$ [29]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [7],\t/a/regfile/regfile$27$ [29]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u379_o,_al_u547_o}),
    .q({\t/a/regfile/regfile$26$ [7],\t/a/regfile/regfile$26$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b840|t/a/regfile/reg0_b853  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [8],\t/a/regfile/regfile$26$ [21]}),
    .e({\t/a/regfile/regfile$27$ [8],\t/a/regfile/regfile$27$ [21]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u372_o,_al_u729_o}),
    .q({\t/a/regfile/regfile$26$ [8],\t/a/regfile/regfile$26$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b841|t/a/regfile/reg0_b859  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$26$ [9],\t/a/regfile/regfile$26$ [27]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [9],\t/a/regfile/regfile$27$ [27]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u337_o,_al_u589_o}),
    .q({\t/a/regfile/regfile$26$ [9],\t/a/regfile/regfile$26$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b842|t/a/regfile/reg0_b851  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [10],\t/a/regfile/regfile$26$ [19]}),
    .e({\t/a/regfile/regfile$27$ [10],\t/a/regfile/regfile$27$ [19]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u981_o,_al_u792_o}),
    .q({\t/a/regfile/regfile$26$ [10],\t/a/regfile/regfile$26$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b843|t/a/regfile/reg0_b854  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$26$ [11],\t/a/regfile/regfile$26$ [22]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [11],\t/a/regfile/regfile$27$ [22]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u946_o,_al_u694_o}),
    .q({\t/a/regfile/regfile$26$ [11],\t/a/regfile/regfile$26$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b844|t/a/regfile/reg0_b849  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [12],\t/a/regfile/regfile$26$ [17]}),
    .e({\t/a/regfile/regfile$27$ [12],\t/a/regfile/regfile$27$ [17]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [17]}),
    .sr(rst_pad),
    .f({_al_u939_o,_al_u834_o}),
    .q({\t/a/regfile/regfile$26$ [12],\t/a/regfile/regfile$26$ [17]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b845|t/a/regfile/reg0_b852  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$26$ [13],\t/a/regfile/regfile$26$ [20]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [13],\t/a/regfile/regfile$27$ [20]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u904_o,_al_u736_o}),
    .q({\t/a/regfile/regfile$26$ [13],\t/a/regfile/regfile$26$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b846|t/a/regfile/reg0_b847  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [14],\t/a/regfile/regfile$26$ [15]}),
    .e({\t/a/regfile/regfile$27$ [14],\t/a/regfile/regfile$27$ [15]}),
    .mi({\t/a/reg_writedat [14],\t/a/reg_writedat [15]}),
    .sr(rst_pad),
    .f({_al_u897_o,_al_u876_o}),
    .q({\t/a/regfile/regfile$26$ [14],\t/a/regfile/regfile$26$ [15]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b848|t/a/regfile/reg0_b850  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$26$ [16],\t/a/regfile/regfile$26$ [18]}),
    .ce(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [16],\t/a/regfile/regfile$27$ [18]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u841_o,_al_u799_o}),
    .q({\t/a/regfile/regfile$26$ [16],\t/a/regfile/regfile$26$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*~D*C*B*A)"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b864|t/a/regfile/reg0_b895  (
    .a({_al_u256_o,\t/a/ID_rs2 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs2 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$26$ [31]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$27$ [31]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b864_sel_is_3_o ,_al_u1214_o}),
    .q({\t/a/regfile/regfile$27$ [0],\t/a/regfile/regfile$27$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b865|t/a/regfile/reg0_b893  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [1],\t/a/regfile/regfile$26$ [29]}),
    .e({\t/a/regfile/regfile$27$ [1],\t/a/regfile/regfile$27$ [29]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u1487_o,_al_u1277_o}),
    .q({\t/a/regfile/regfile$27$ [1],\t/a/regfile/regfile$27$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b866|t/a/regfile/reg0_b891  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [2],\t/a/regfile/regfile$26$ [27]}),
    .e({\t/a/regfile/regfile$27$ [2],\t/a/regfile/regfile$27$ [27]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u1256_o,_al_u1319_o}),
    .q({\t/a/regfile/regfile$27$ [2],\t/a/regfile/regfile$27$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000010010001100),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000010010001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b867|t/a/regfile/reg0_b878  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$26$ [3],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [3],\t/a/regfile/regfile$26$ [14]}),
    .e({open_n29032,\t/a/regfile/regfile$27$ [14]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [14]}),
    .sr(rst_pad),
    .f({_al_u1179_o,_al_u1613_o}),
    .q({\t/a/regfile/regfile$27$ [3],\t/a/regfile/regfile$27$ [14]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b868|t/a/regfile/reg0_b889  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [4],\t/a/regfile/regfile$26$ [25]}),
    .e({\t/a/regfile/regfile$27$ [4],\t/a/regfile/regfile$27$ [25]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [25]}),
    .sr(rst_pad),
    .f({_al_u1172_o,_al_u1361_o}),
    .q({\t/a/regfile/regfile$27$ [4],\t/a/regfile/regfile$27$ [25]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b869|t/a/regfile/reg0_b888  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [5],\t/a/regfile/regfile$26$ [24]}),
    .e({\t/a/regfile/regfile$27$ [5],\t/a/regfile/regfile$27$ [24]}),
    .mi({\t/a/reg_writedat [5],\t/a/reg_writedat [24]}),
    .sr(rst_pad),
    .f({_al_u1151_o,_al_u1382_o}),
    .q({\t/a/regfile/regfile$27$ [5],\t/a/regfile/regfile$27$ [24]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b870|t/a/regfile/reg0_b886  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [6],\t/a/regfile/regfile$26$ [22]}),
    .e({\t/a/regfile/regfile$27$ [6],\t/a/regfile/regfile$27$ [22]}),
    .mi({\t/a/reg_writedat [6],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u1130_o,_al_u1424_o}),
    .q({\t/a/regfile/regfile$27$ [6],\t/a/regfile/regfile$27$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b871|t/a/regfile/reg0_b884  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [7],\t/a/regfile/regfile$26$ [20]}),
    .e({\t/a/regfile/regfile$27$ [7],\t/a/regfile/regfile$27$ [20]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u1109_o,_al_u1466_o}),
    .q({\t/a/regfile/regfile$27$ [7],\t/a/regfile/regfile$27$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b872|t/a/regfile/reg0_b894  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$26$ [8],\t/a/regfile/regfile$26$ [30]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [8],\t/a/regfile/regfile$27$ [30]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1074_o,_al_u1221_o}),
    .q({\t/a/regfile/regfile$27$ [8],\t/a/regfile/regfile$27$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b873|t/a/regfile/reg0_b883  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [9],\t/a/regfile/regfile$26$ [19]}),
    .e({\t/a/regfile/regfile$27$ [9],\t/a/regfile/regfile$27$ [19]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [19]}),
    .sr(rst_pad),
    .f({_al_u1067_o,_al_u1508_o}),
    .q({\t/a/regfile/regfile$27$ [9],\t/a/regfile/regfile$27$ [19]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b874|t/a/regfile/reg0_b892  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$26$ [10],\t/a/regfile/regfile$26$ [28]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [10],\t/a/regfile/regfile$27$ [28]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1683_o,_al_u1284_o}),
    .q({\t/a/regfile/regfile$27$ [10],\t/a/regfile/regfile$27$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b875|t/a/regfile/reg0_b882  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [11],\t/a/regfile/regfile$26$ [18]}),
    .e({\t/a/regfile/regfile$27$ [11],\t/a/regfile/regfile$27$ [18]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u1676_o,_al_u1529_o}),
    .q({\t/a/regfile/regfile$27$ [11],\t/a/regfile/regfile$27$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b876|t/a/regfile/reg0_b890  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$26$ [12],\t/a/regfile/regfile$26$ [26]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [12],\t/a/regfile/regfile$27$ [26]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1641_o,_al_u1326_o}),
    .q({\t/a/regfile/regfile$27$ [12],\t/a/regfile/regfile$27$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(~C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(~C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000011100000011),
    .INIT_LUTF1(16'b0000011100000011),
    .INIT_LUTG0(16'b0000111100001011),
    .INIT_LUTG1(16'b0000111100001011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b877|t/a/regfile/reg0_b880  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$26$ [13],\t/a/regfile/regfile$26$ [16]}),
    .e({\t/a/regfile/regfile$27$ [13],\t/a/regfile/regfile$27$ [16]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [16]}),
    .sr(rst_pad),
    .f({_al_u1634_o,_al_u1571_o}),
    .q({\t/a/regfile/regfile$27$ [13],\t/a/regfile/regfile$27$ [16]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b879|t/a/regfile/reg0_b887  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$26$ [15],\t/a/regfile/regfile$26$ [23]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [15],\t/a/regfile/regfile$27$ [23]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1578_o,_al_u1389_o}),
    .q({\t/a/regfile/regfile$27$ [15],\t/a/regfile/regfile$27$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000010010001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b881|t/a/regfile/reg0_b885  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$26$ [17],\t/a/regfile/regfile$26$ [21]}),
    .ce(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$27$ [17],\t/a/regfile/regfile$27$ [21]}),
    .mi({\t/a/reg_writedat [17],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1536_o,_al_u1431_o}),
    .q({\t/a/regfile/regfile$27$ [17],\t/a/regfile/regfile$27$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b900|t/a/regfile/reg0_b927  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$28$ [4],\t/a/regfile/regfile$28$ [31]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [4],\t/a/regfile/regfile$29$ [31]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u439_o,_al_u481_o}),
    .q({\t/a/regfile/regfile$28$ [4],\t/a/regfile/regfile$28$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b903|t/a/regfile/reg0_b925  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$28$ [7],\t/a/regfile/regfile$28$ [29]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [7],\t/a/regfile/regfile$29$ [29]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u376_o,_al_u544_o}),
    .q({\t/a/regfile/regfile$28$ [7],\t/a/regfile/regfile$28$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b905|t/a/regfile/reg0_b923  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$28$ [9],\t/a/regfile/regfile$28$ [27]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [9],\t/a/regfile/regfile$29$ [27]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u334_o,_al_u586_o}),
    .q({\t/a/regfile/regfile$28$ [9],\t/a/regfile/regfile$28$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b907|t/a/regfile/reg0_b918  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$28$ [11],\t/a/regfile/regfile$28$ [22]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [11],\t/a/regfile/regfile$29$ [22]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u943_o,_al_u691_o}),
    .q({\t/a/regfile/regfile$28$ [11],\t/a/regfile/regfile$28$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b909|t/a/regfile/reg0_b916  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$28$ [13],\t/a/regfile/regfile$28$ [20]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [13],\t/a/regfile/regfile$29$ [20]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u901_o,_al_u733_o}),
    .q({\t/a/regfile/regfile$28$ [13],\t/a/regfile/regfile$28$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b912|t/a/regfile/reg0_b914  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$28$ [16],\t/a/regfile/regfile$28$ [18]}),
    .ce(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [16],\t/a/regfile/regfile$29$ [18]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u838_o,_al_u796_o}),
    .q({\t/a/regfile/regfile$28$ [16],\t/a/regfile/regfile$28$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b931|t/a/regfile/reg0_b958  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$28$ [3],\t/a/regfile/regfile$28$ [30]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [3],\t/a/regfile/regfile$29$ [30]}),
    .mi({\t/a/reg_writedat [3],\t/a/reg_writedat [30]}),
    .sr(rst_pad),
    .f({_al_u1176_o,_al_u1218_o}),
    .q({\t/a/regfile/regfile$29$ [3],\t/a/regfile/regfile$29$ [30]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b936|t/a/regfile/reg0_b956  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$28$ [8],\t/a/regfile/regfile$28$ [28]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [8],\t/a/regfile/regfile$29$ [28]}),
    .mi({\t/a/reg_writedat [8],\t/a/reg_writedat [28]}),
    .sr(rst_pad),
    .f({_al_u1071_o,_al_u1281_o}),
    .q({\t/a/regfile/regfile$29$ [8],\t/a/regfile/regfile$29$ [28]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b938|t/a/regfile/reg0_b954  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$28$ [10],\t/a/regfile/regfile$28$ [26]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [10],\t/a/regfile/regfile$29$ [26]}),
    .mi({\t/a/reg_writedat [10],\t/a/reg_writedat [26]}),
    .sr(rst_pad),
    .f({_al_u1680_o,_al_u1323_o}),
    .q({\t/a/regfile/regfile$29$ [10],\t/a/regfile/regfile$29$ [26]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b940|t/a/regfile/reg0_b951  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$28$ [12],\t/a/regfile/regfile$28$ [23]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [12],\t/a/regfile/regfile$29$ [23]}),
    .mi({\t/a/reg_writedat [12],\t/a/reg_writedat [23]}),
    .sr(rst_pad),
    .f({_al_u1638_o,_al_u1386_o}),
    .q({\t/a/regfile/regfile$29$ [12],\t/a/regfile/regfile$29$ [23]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    //.LUT1("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100100011),
    .INIT_LUT1(16'b0000000100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b943|t/a/regfile/reg0_b949  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/regfile/regfile$28$ [15],\t/a/regfile/regfile$28$ [21]}),
    .ce(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$29$ [15],\t/a/regfile/regfile$29$ [21]}),
    .mi({\t/a/reg_writedat [15],\t/a/reg_writedat [21]}),
    .sr(rst_pad),
    .f({_al_u1575_o,_al_u1428_o}),
    .q({\t/a/regfile/regfile$29$ [15],\t/a/regfile/regfile$29$ [21]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(0*D*C*~B*A)"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(1*D*C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b960|t/a/regfile/reg0_b966  (
    .a({_al_u256_o,\t/a/ID_rs1 [0]}),
    .b({\t/a/WB_rd [0],\t/a/ID_rs1 [1]}),
    .c({\t/a/WB_rd [1],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/WB_rd [2],\t/a/regfile/regfile$30$ [6]}),
    .e({\t/a/WB_rd [3],\t/a/regfile/regfile$31$ [6]}),
    .mi({\t/a/reg_writedat [0],\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({\t/a/regfile/mux39_b960_sel_is_3_o ,_al_u412_o}),
    .q({\t/a/regfile/regfile$30$ [0],\t/a/regfile/regfile$30$ [6]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b961|t/a/regfile/reg0_b965  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [1],\t/a/regfile/regfile$30$ [5]}),
    .e({\t/a/regfile/regfile$31$ [1],\t/a/regfile/regfile$31$ [5]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u769_o,_al_u433_o}),
    .q({\t/a/regfile/regfile$30$ [1],\t/a/regfile/regfile$30$ [5]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b962|t/a/regfile/reg0_b963  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/ID_rs1 [2],\t/a/ID_rs1 [2]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [2],\t/a/regfile/regfile$30$ [3]}),
    .e({\t/a/regfile/regfile$31$ [2],\t/a/regfile/regfile$31$ [3]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [3]}),
    .sr(rst_pad),
    .f({_al_u538_o,_al_u475_o}),
    .q({\t/a/regfile/regfile$30$ [2],\t/a/regfile/regfile$30$ [3]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b964|t/a/regfile/reg0_b991  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$30$ [4],\t/a/regfile/regfile$31$ [31]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$31$ [4],\t/a/regfile/regfile$30$ [31]}),
    .mi({\t/a/reg_writedat [4],\t/a/reg_writedat [31]}),
    .sr(rst_pad),
    .f({_al_u440_o,_al_u482_o}),
    .q({\t/a/regfile/regfile$30$ [4],\t/a/regfile/regfile$30$ [31]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000010010001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b967|t/a/regfile/reg0_b989  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$30$ [7],\t/a/regfile/regfile$31$ [29]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$31$ [7],\t/a/regfile/regfile$30$ [29]}),
    .mi({\t/a/reg_writedat [7],\t/a/reg_writedat [29]}),
    .sr(rst_pad),
    .f({_al_u377_o,_al_u545_o}),
    .q({\t/a/regfile/regfile$30$ [7],\t/a/regfile/regfile$30$ [29]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b969|t/a/regfile/reg0_b987  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [9],\t/a/regfile/regfile$31$ [27]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [9],\t/a/regfile/regfile$30$ [27]}),
    .mi({\t/a/reg_writedat [9],\t/a/reg_writedat [27]}),
    .sr(rst_pad),
    .f({_al_u335_o,_al_u587_o}),
    .q({\t/a/regfile/regfile$30$ [9],\t/a/regfile/regfile$30$ [27]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b971|t/a/regfile/reg0_b982  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [11],\t/a/regfile/regfile$31$ [22]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [11],\t/a/regfile/regfile$30$ [22]}),
    .mi({\t/a/reg_writedat [11],\t/a/reg_writedat [22]}),
    .sr(rst_pad),
    .f({_al_u944_o,_al_u692_o}),
    .q({\t/a/regfile/regfile$30$ [11],\t/a/regfile/regfile$30$ [22]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b973|t/a/regfile/reg0_b980  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [13],\t/a/regfile/regfile$31$ [20]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [13],\t/a/regfile/regfile$30$ [20]}),
    .mi({\t/a/reg_writedat [13],\t/a/reg_writedat [20]}),
    .sr(rst_pad),
    .f({_al_u902_o,_al_u734_o}),
    .q({\t/a/regfile/regfile$30$ [13],\t/a/regfile/regfile$30$ [20]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_MSLICE #(
    //.LUT0("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    //.LUT1("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100001001100),
    .INIT_LUT1(16'b0000100001001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b976|t/a/regfile/reg0_b978  (
    .a({\t/a/ID_rs1 [0],\t/a/ID_rs1 [0]}),
    .b({\t/a/ID_rs1 [1],\t/a/ID_rs1 [1]}),
    .c({\t/a/regfile/regfile$31$ [16],\t/a/regfile/regfile$31$ [18]}),
    .ce(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [16],\t/a/regfile/regfile$30$ [18]}),
    .mi({\t/a/reg_writedat [16],\t/a/reg_writedat [18]}),
    .sr(rst_pad),
    .f({_al_u839_o,_al_u797_o}),
    .q({\t/a/regfile/regfile$30$ [16],\t/a/regfile/regfile$30$ [18]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b993|t/a/regfile/reg0_b998  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [1],\t/a/regfile/regfile$30$ [6]}),
    .e({\t/a/regfile/regfile$31$ [1],\t/a/regfile/regfile$31$ [6]}),
    .mi({\t/a/reg_writedat [1],\t/a/reg_writedat [6]}),
    .sr(rst_pad),
    .f({_al_u1485_o,_al_u1128_o}),
    .q({\t/a/regfile/regfile$31$ [1],\t/a/regfile/regfile$31$ [6]}));  // register.v(63)
  // register.v(63)
  // register.v(63)
  EG_PHY_LSLICE #(
    //.LUTF0("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTF1("(C*~(B*~(D*~(0)*~(A)+D*0*~(A)+~(D)*0*A+D*0*A)))"),
    //.LUTG0("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    //.LUTG1("(C*~(B*~(D*~(1)*~(A)+D*1*~(A)+~(D)*1*A+D*1*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111000000110000),
    .INIT_LUTF1(16'b0111000000110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("MI"),
    .REG1_REGSET("SET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \t/a/regfile/reg0_b994|t/a/regfile/reg0_b997  (
    .a({\t/a/ID_rs2 [0],\t/a/ID_rs2 [0]}),
    .b({\t/a/ID_rs2 [1],\t/a/ID_rs2 [1]}),
    .c({\t/a/ID_rs2 [2],\t/a/ID_rs2 [2]}),
    .ce(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .clk(clock_pad),
    .d({\t/a/regfile/regfile$30$ [2],\t/a/regfile/regfile$30$ [5]}),
    .e({\t/a/regfile/regfile$31$ [2],\t/a/regfile/regfile$31$ [5]}),
    .mi({\t/a/reg_writedat [2],\t/a/reg_writedat [5]}),
    .sr(rst_pad),
    .f({_al_u1254_o,_al_u1149_o}),
    .q({\t/a/regfile/regfile$31$ [2],\t/a/regfile/regfile$31$ [5]}));  // register.v(63)
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u1/u0|u1/ucin  (
    .a({\t/memstraddress [2],1'b0}),
    .b({1'b1,open_n29514}),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .mi({open_n29529,\t/memstraddress [2]}),
    .sr(rst_pad),
    .f({n4[0],open_n29530}),
    .fco(\u1/c1 ),
    .q({open_n29533,\t/a/ID_memstraddr [2]}));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u10|u1/u9  (
    .a(\t/memstraddress [12:11]),
    .b(2'b00),
    .fci(\u1/c9 ),
    .f(n4[10:9]),
    .fco(\u1/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u12|u1/u11  (
    .a(\t/memstraddress [14:13]),
    .b(2'b00),
    .fci(\u1/c11 ),
    .f(n4[12:11]),
    .fco(\u1/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u14|u1/u13  (
    .a(\t/memstraddress [16:15]),
    .b(2'b00),
    .fci(\u1/c13 ),
    .f(n4[14:13]),
    .fco(\u1/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u16|u1/u15  (
    .a(\t/memstraddress [18:17]),
    .b(2'b00),
    .fci(\u1/c15 ),
    .f(n4[16:15]),
    .fco(\u1/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u18|u1/u17  (
    .a(\t/memstraddress [20:19]),
    .b(2'b00),
    .fci(\u1/c17 ),
    .f(n4[18:17]),
    .fco(\u1/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u20|u1/u19  (
    .a(\t/memstraddress [22:21]),
    .b(2'b00),
    .fci(\u1/c19 ),
    .f(n4[20:19]),
    .fco(\u1/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u22|u1/u21  (
    .a(\t/memstraddress [24:23]),
    .b(2'b00),
    .fci(\u1/c21 ),
    .f(n4[22:21]),
    .fco(\u1/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u24|u1/u23  (
    .a(\t/memstraddress [26:25]),
    .b(2'b00),
    .fci(\u1/c23 ),
    .f(n4[24:23]),
    .fco(\u1/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u26|u1/u25  (
    .a(\t/memstraddress [28:27]),
    .b(2'b00),
    .fci(\u1/c25 ),
    .f(n4[26:25]),
    .fco(\u1/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u28|u1/u27  (
    .a(\t/memstraddress [30:29]),
    .b(2'b00),
    .fci(\u1/c27 ),
    .f(n4[28:27]),
    .fco(\u1/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u29_al_u2978  (
    .a({open_n29754,\t/memstraddress [31]}),
    .b({open_n29755,1'b0}),
    .fci(\u1/c29 ),
    .f({open_n29774,n4[29]}));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u2|u1/u1  (
    .a(\t/memstraddress [4:3]),
    .b(2'b00),
    .fci(\u1/c1 ),
    .f(n4[2:1]),
    .fco(\u1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u4|u1/u3  (
    .a(\t/memstraddress [6:5]),
    .b(2'b00),
    .fci(\u1/c3 ),
    .f(n4[4:3]),
    .fco(\u1/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u6|u1/u5  (
    .a(\t/memstraddress [8:7]),
    .b(2'b00),
    .fci(\u1/c5 ),
    .f(n4[6:5]),
    .fco(\u1/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u1/u8|u1/u7  (
    .a(\t/memstraddress [10:9]),
    .b(2'b00),
    .fci(\u1/c7 ),
    .f(n4[8:7]),
    .fco(\u1/c9 ));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u11_al_u2964  (
    .a({\t/a/ID_jump_addr [14],\t/a/ID_jump_addr [12]}),
    .b({\t/a/ID_jump_addr [15],\t/a/ID_jump_addr [13]}),
    .c(2'b00),
    .d({n4[12],n4[10]}),
    .e({n4[13],n4[11]}),
    .fci(\u3/c11 ),
    .f({n8[13],n8[11]}),
    .fco(\u3/c15 ),
    .fx({n8[14],n8[12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u15_al_u2965  (
    .a({\t/a/ID_jump_addr [18],\t/a/ID_jump_addr [16]}),
    .b({\t/a/ID_jump_addr [19],\t/a/ID_jump_addr [17]}),
    .c(2'b00),
    .d({n4[16],n4[14]}),
    .e({n4[17],n4[15]}),
    .fci(\u3/c15 ),
    .f({n8[17],n8[15]}),
    .fco(\u3/c19 ),
    .fx({n8[18],n8[16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u19_al_u2966  (
    .a({\t/a/ID_jump_addr [22],\t/a/ID_jump_addr [20]}),
    .b({\t/a/ID_jump_addr [23],\t/a/ID_jump_addr [21]}),
    .c(2'b00),
    .d({n4[20],n4[18]}),
    .e({n4[21],n4[19]}),
    .fci(\u3/c19 ),
    .f({n8[21],n8[19]}),
    .fco(\u3/c23 ),
    .fx({n8[22],n8[20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u23_al_u2967  (
    .a({\t/a/ID_jump_addr [26],\t/a/ID_jump_addr [24]}),
    .b({\t/a/ID_jump_addr [27],\t/a/ID_jump_addr [25]}),
    .c(2'b00),
    .d({n4[24],n4[22]}),
    .e({n4[25],n4[23]}),
    .fci(\u3/c23 ),
    .f({n8[25],n8[23]}),
    .fco(\u3/c27 ),
    .fx({n8[26],n8[24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u27_al_u2968  (
    .a({\t/a/ID_jump_addr [30],\t/a/ID_jump_addr [28]}),
    .b({\t/a/ID_jump_addr [31],\t/a/ID_jump_addr [29]}),
    .c(2'b00),
    .d({n4[28],n4[26]}),
    .e({n4[29],n4[27]}),
    .fci(\u3/c27 ),
    .f({n8[29],n8[27]}),
    .fx({n8[30],n8[28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u3_al_u2962  (
    .a({\t/a/ID_jump_addr [6],\t/a/ID_jump_addr [4]}),
    .b({\t/a/ID_jump_addr [7],\t/a/ID_jump_addr [5]}),
    .c(2'b00),
    .d({n4[4],n4[2]}),
    .e({n4[5],n4[3]}),
    .fci(\u3/c3 ),
    .f({n8[5],n8[3]}),
    .fco(\u3/c7 ),
    .fx({n8[6],n8[4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u3/u7_al_u2963  (
    .a({\t/a/ID_jump_addr [10],\t/a/ID_jump_addr [8]}),
    .b({\t/a/ID_jump_addr [11],\t/a/ID_jump_addr [9]}),
    .c(2'b00),
    .d({n4[8],n4[6]}),
    .e({n4[9],n4[7]}),
    .fci(\u3/c7 ),
    .f({n8[9],n8[7]}),
    .fco(\u3/c11 ),
    .fx({n8[10],n8[8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u3/ucin_al_u2961"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u3/ucin_al_u2961  (
    .a({\t/a/ID_jump_addr [2],1'b0}),
    .b({\t/a/ID_jump_addr [3],\t/a/ID_jump_addr [1]}),
    .c(2'b00),
    .ce(\t/a/if_id/n9 ),
    .clk(clock_pad),
    .d({n4[0],1'b1}),
    .e({n4[1],\t/memstraddress [1]}),
    .mi({open_n29996,\t/memstraddress [1]}),
    .sr(rst_pad),
    .f({n8[1],open_n30008}),
    .fco(\u3/c3 ),
    .fx({n8[2],n8[0]}),
    .q({open_n30009,\t/a/ID_memstraddr [1]}));

endmodule 

