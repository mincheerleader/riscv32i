// Verilog netlist created by TD v4.3.815
// Fri Mar 22 13:53:33 2019

`timescale 1ns / 1ps
module __top  // __top.v(3)
  (
  clock,
  rst,
  led
  );

  input clock;  // __top.v(4)
  input rst;  // __top.v(3)
  output led;  // __top.v(5)

  wire [31:0] addr;  // __top.v(17)
  wire [31:0] i_data;  // __top.v(15)
  wire [3:0] n2;
  wire [3:0] n3;
  wire [31:0] o_data;  // __top.v(16)
  wire [31:0] \t/a/EX_A ;  // cpu.v(47)
  wire [31:0] \t/a/EX_B ;  // cpu.v(48)
  wire [2:0] \t/a/EX_fun3 ;  // cpu.v(49)
  wire [6:0] \t/a/EX_fun7 ;  // cpu.v(41)
  wire [31:0] \t/a/EX_memstraddr ;  // cpu.v(38)
  wire [6:0] \t/a/EX_op ;  // cpu.v(42)
  wire [3:0] \t/a/EX_operation ;  // cpu.v(46)
  wire [4:0] \t/a/EX_rd ;  // cpu.v(45)
  wire [31:0] \t/a/EX_regdat1 ;  // cpu.v(39)
  wire [31:0] \t/a/EX_regdat2 ;  // cpu.v(40)
  wire [4:0] \t/a/EX_rs1 ;  // cpu.v(43)
  wire [4:0] \t/a/EX_rs2 ;  // cpu.v(44)
  wire [2:0] \t/a/ID_fun3 ;  // cpu.v(21)
  wire [6:0] \t/a/ID_fun7 ;  // cpu.v(22)
  wire [31:0] \t/a/ID_jump_addr ;  // cpu.v(28)
  wire [31:0] \t/a/ID_jump_regdat1 ;  // cpu.v(29)
  wire [31:0] \t/a/ID_jump_regdat2 ;  // cpu.v(30)
  wire [31:0] \t/a/ID_memstraddr ;  // cpu.v(26)
  wire [6:0] \t/a/ID_op ;  // cpu.v(20)
  wire [4:0] \t/a/ID_rd ;  // cpu.v(23)
  wire [31:0] \t/a/ID_read_dat1 ;  // cpu.v(36)
  wire [31:0] \t/a/ID_read_dat2 ;  // cpu.v(37)
  wire [4:0] \t/a/ID_rs1 ;  // cpu.v(24)
  wire [4:0] \t/a/ID_rs2 ;  // cpu.v(25)
  wire [31:0] \t/a/IF_skip_addr ;  // cpu.v(17)
  wire [31:0] \t/a/MEM_aludat ;  // cpu.v(54)
  wire [2:0] \t/a/MEM_fun3 ;  // cpu.v(58)
  wire [6:0] \t/a/MEM_op ;  // cpu.v(55)
  wire [4:0] \t/a/MEM_rd ;  // cpu.v(56)
  wire [31:0] \t/a/MEM_regdat2 ;  // cpu.v(57)
  wire [6:0] \t/a/WB_op ;  // cpu.v(71)
  wire [4:0] \t/a/WB_rd ;  // cpu.v(70)
  wire [31:0] \t/a/alu/n12 ;
  wire [31:0] \t/a/alu/n14 ;
  wire [31:0] \t/a/alu/n15 ;
  wire [31:0] \t/a/alu/n48 ;
  wire [31:0] \t/a/alu/n49 ;
  wire [31:0] \t/a/alu/n5 ;
  wire [31:0] \t/a/alu/n6 ;
  wire [31:0] \t/a/alu/n7 ;
  wire [1:0] \t/a/alu_A_select ;  // cpu.v(33)
  wire [1:0] \t/a/alu_B_select ;  // cpu.v(34)
  wire [31:0] \t/a/aludat ;  // cpu.v(52)
  wire [3:0] \t/a/aluin/n40 ;
  wire [3:0] \t/a/aluin/n41 ;
  wire [6:0] \t/a/aluin/n9 ;
  wire [31:0] \t/a/aluin/o_A1 ;  // alu.v(25)
  wire [31:0] \t/a/aluin/o_B1 ;  // alu.v(24)
  wire [3:0] \t/a/aluin/operation_R ;  // alu.v(22)
  wire  \t/a/aluin/sel0_b0/B0 ;
  wire  \t/a/aluin/sel0_b0/B1 ;
  wire  \t/a/aluin/sel0_b0/B2 ;
  wire  \t/a/aluin/sel0_b0/B3 ;
  wire  \t/a/aluin/sel0_b1/B0 ;
  wire  \t/a/aluin/sel0_b1/B1 ;
  wire  \t/a/aluin/sel0_b1/B2 ;
  wire  \t/a/aluin/sel0_b1/B3 ;
  wire  \t/a/aluin/sel0_b10/B0 ;
  wire  \t/a/aluin/sel0_b10/B1 ;
  wire  \t/a/aluin/sel0_b10/B2 ;
  wire  \t/a/aluin/sel0_b10/B3 ;
  wire  \t/a/aluin/sel0_b11/B0 ;
  wire  \t/a/aluin/sel0_b11/B1 ;
  wire  \t/a/aluin/sel0_b11/B2 ;
  wire  \t/a/aluin/sel0_b11/B3 ;
  wire  \t/a/aluin/sel0_b12/B0 ;
  wire  \t/a/aluin/sel0_b12/B1 ;
  wire  \t/a/aluin/sel0_b12/B2 ;
  wire  \t/a/aluin/sel0_b12/B3 ;
  wire  \t/a/aluin/sel0_b13/B0 ;
  wire  \t/a/aluin/sel0_b13/B1 ;
  wire  \t/a/aluin/sel0_b13/B2 ;
  wire  \t/a/aluin/sel0_b13/B3 ;
  wire  \t/a/aluin/sel0_b14/B0 ;
  wire  \t/a/aluin/sel0_b14/B1 ;
  wire  \t/a/aluin/sel0_b14/B2 ;
  wire  \t/a/aluin/sel0_b14/B3 ;
  wire  \t/a/aluin/sel0_b15/B0 ;
  wire  \t/a/aluin/sel0_b15/B1 ;
  wire  \t/a/aluin/sel0_b15/B2 ;
  wire  \t/a/aluin/sel0_b15/B3 ;
  wire  \t/a/aluin/sel0_b16/B0 ;
  wire  \t/a/aluin/sel0_b16/B1 ;
  wire  \t/a/aluin/sel0_b16/B2 ;
  wire  \t/a/aluin/sel0_b16/B3 ;
  wire  \t/a/aluin/sel0_b17/B0 ;
  wire  \t/a/aluin/sel0_b17/B1 ;
  wire  \t/a/aluin/sel0_b17/B2 ;
  wire  \t/a/aluin/sel0_b17/B3 ;
  wire  \t/a/aluin/sel0_b18/B0 ;
  wire  \t/a/aluin/sel0_b18/B1 ;
  wire  \t/a/aluin/sel0_b18/B2 ;
  wire  \t/a/aluin/sel0_b18/B3 ;
  wire  \t/a/aluin/sel0_b19/B0 ;
  wire  \t/a/aluin/sel0_b19/B1 ;
  wire  \t/a/aluin/sel0_b19/B2 ;
  wire  \t/a/aluin/sel0_b19/B3 ;
  wire  \t/a/aluin/sel0_b2/B0 ;
  wire  \t/a/aluin/sel0_b2/B1 ;
  wire  \t/a/aluin/sel0_b2/B2 ;
  wire  \t/a/aluin/sel0_b2/B3 ;
  wire  \t/a/aluin/sel0_b20/B0 ;
  wire  \t/a/aluin/sel0_b20/B1 ;
  wire  \t/a/aluin/sel0_b20/B2 ;
  wire  \t/a/aluin/sel0_b20/B3 ;
  wire  \t/a/aluin/sel0_b21/B0 ;
  wire  \t/a/aluin/sel0_b21/B1 ;
  wire  \t/a/aluin/sel0_b21/B2 ;
  wire  \t/a/aluin/sel0_b21/B3 ;
  wire  \t/a/aluin/sel0_b22/B0 ;
  wire  \t/a/aluin/sel0_b22/B1 ;
  wire  \t/a/aluin/sel0_b22/B2 ;
  wire  \t/a/aluin/sel0_b22/B3 ;
  wire  \t/a/aluin/sel0_b23/B0 ;
  wire  \t/a/aluin/sel0_b23/B1 ;
  wire  \t/a/aluin/sel0_b23/B2 ;
  wire  \t/a/aluin/sel0_b23/B3 ;
  wire  \t/a/aluin/sel0_b24/B0 ;
  wire  \t/a/aluin/sel0_b24/B1 ;
  wire  \t/a/aluin/sel0_b24/B2 ;
  wire  \t/a/aluin/sel0_b24/B3 ;
  wire  \t/a/aluin/sel0_b25/B0 ;
  wire  \t/a/aluin/sel0_b25/B1 ;
  wire  \t/a/aluin/sel0_b25/B2 ;
  wire  \t/a/aluin/sel0_b25/B3 ;
  wire  \t/a/aluin/sel0_b26/B0 ;
  wire  \t/a/aluin/sel0_b26/B1 ;
  wire  \t/a/aluin/sel0_b26/B2 ;
  wire  \t/a/aluin/sel0_b26/B3 ;
  wire  \t/a/aluin/sel0_b27/B0 ;
  wire  \t/a/aluin/sel0_b27/B1 ;
  wire  \t/a/aluin/sel0_b27/B2 ;
  wire  \t/a/aluin/sel0_b27/B3 ;
  wire  \t/a/aluin/sel0_b28/B0 ;
  wire  \t/a/aluin/sel0_b28/B1 ;
  wire  \t/a/aluin/sel0_b28/B2 ;
  wire  \t/a/aluin/sel0_b28/B3 ;
  wire  \t/a/aluin/sel0_b29/B0 ;
  wire  \t/a/aluin/sel0_b29/B1 ;
  wire  \t/a/aluin/sel0_b29/B2 ;
  wire  \t/a/aluin/sel0_b29/B3 ;
  wire  \t/a/aluin/sel0_b3/B0 ;
  wire  \t/a/aluin/sel0_b3/B1 ;
  wire  \t/a/aluin/sel0_b3/B2 ;
  wire  \t/a/aluin/sel0_b3/B3 ;
  wire  \t/a/aluin/sel0_b30/B0 ;
  wire  \t/a/aluin/sel0_b30/B1 ;
  wire  \t/a/aluin/sel0_b30/B2 ;
  wire  \t/a/aluin/sel0_b30/B3 ;
  wire  \t/a/aluin/sel0_b31/B0 ;
  wire  \t/a/aluin/sel0_b31/B1 ;
  wire  \t/a/aluin/sel0_b31/B2 ;
  wire  \t/a/aluin/sel0_b31/B3 ;
  wire  \t/a/aluin/sel0_b4/B0 ;
  wire  \t/a/aluin/sel0_b4/B1 ;
  wire  \t/a/aluin/sel0_b4/B2 ;
  wire  \t/a/aluin/sel0_b4/B3 ;
  wire  \t/a/aluin/sel0_b5/B0 ;
  wire  \t/a/aluin/sel0_b5/B1 ;
  wire  \t/a/aluin/sel0_b5/B2 ;
  wire  \t/a/aluin/sel0_b5/B3 ;
  wire  \t/a/aluin/sel0_b6/B0 ;
  wire  \t/a/aluin/sel0_b6/B1 ;
  wire  \t/a/aluin/sel0_b6/B2 ;
  wire  \t/a/aluin/sel0_b6/B3 ;
  wire  \t/a/aluin/sel0_b7/B0 ;
  wire  \t/a/aluin/sel0_b7/B1 ;
  wire  \t/a/aluin/sel0_b7/B2 ;
  wire  \t/a/aluin/sel0_b7/B3 ;
  wire  \t/a/aluin/sel0_b8/B0 ;
  wire  \t/a/aluin/sel0_b8/B1 ;
  wire  \t/a/aluin/sel0_b8/B2 ;
  wire  \t/a/aluin/sel0_b8/B3 ;
  wire  \t/a/aluin/sel0_b9/B0 ;
  wire  \t/a/aluin/sel0_b9/B1 ;
  wire  \t/a/aluin/sel0_b9/B2 ;
  wire  \t/a/aluin/sel0_b9/B3 ;
  wire  \t/a/aluin/sel1_b0/B6 ;
  wire  \t/a/aluin/sel1_b0/B7 ;
  wire  \t/a/aluin/sel1_b0/B8 ;
  wire  \t/a/aluin/sel1_b0/B9 ;
  wire  \t/a/aluin/sel1_b1/B6 ;
  wire  \t/a/aluin/sel1_b1/B7 ;
  wire  \t/a/aluin/sel1_b1/B8 ;
  wire  \t/a/aluin/sel1_b1/B9 ;
  wire  \t/a/aluin/sel1_b10/B6 ;
  wire  \t/a/aluin/sel1_b10/B7 ;
  wire  \t/a/aluin/sel1_b10/B8 ;
  wire  \t/a/aluin/sel1_b10/B9 ;
  wire  \t/a/aluin/sel1_b11/B6 ;
  wire  \t/a/aluin/sel1_b11/B7 ;
  wire  \t/a/aluin/sel1_b11/B8 ;
  wire  \t/a/aluin/sel1_b11/B9 ;
  wire  \t/a/aluin/sel1_b12/B2 ;
  wire  \t/a/aluin/sel1_b12/B3 ;
  wire  \t/a/aluin/sel1_b12/B9 ;
  wire  \t/a/aluin/sel1_b13/B2 ;
  wire  \t/a/aluin/sel1_b13/B3 ;
  wire  \t/a/aluin/sel1_b13/B9 ;
  wire  \t/a/aluin/sel1_b14/B2 ;
  wire  \t/a/aluin/sel1_b14/B3 ;
  wire  \t/a/aluin/sel1_b14/B9 ;
  wire  \t/a/aluin/sel1_b15/B2 ;
  wire  \t/a/aluin/sel1_b15/B3 ;
  wire  \t/a/aluin/sel1_b15/B9 ;
  wire  \t/a/aluin/sel1_b16/B2 ;
  wire  \t/a/aluin/sel1_b16/B3 ;
  wire  \t/a/aluin/sel1_b16/B9 ;
  wire  \t/a/aluin/sel1_b17/B2 ;
  wire  \t/a/aluin/sel1_b17/B3 ;
  wire  \t/a/aluin/sel1_b17/B9 ;
  wire  \t/a/aluin/sel1_b18/B2 ;
  wire  \t/a/aluin/sel1_b18/B3 ;
  wire  \t/a/aluin/sel1_b18/B9 ;
  wire  \t/a/aluin/sel1_b19/B2 ;
  wire  \t/a/aluin/sel1_b19/B3 ;
  wire  \t/a/aluin/sel1_b19/B9 ;
  wire  \t/a/aluin/sel1_b2/B6 ;
  wire  \t/a/aluin/sel1_b2/B7 ;
  wire  \t/a/aluin/sel1_b2/B8 ;
  wire  \t/a/aluin/sel1_b2/B9 ;
  wire  \t/a/aluin/sel1_b20/B2 ;
  wire  \t/a/aluin/sel1_b20/B3 ;
  wire  \t/a/aluin/sel1_b20/B9 ;
  wire  \t/a/aluin/sel1_b21/B2 ;
  wire  \t/a/aluin/sel1_b21/B3 ;
  wire  \t/a/aluin/sel1_b21/B9 ;
  wire  \t/a/aluin/sel1_b22/B2 ;
  wire  \t/a/aluin/sel1_b22/B3 ;
  wire  \t/a/aluin/sel1_b22/B9 ;
  wire  \t/a/aluin/sel1_b23/B2 ;
  wire  \t/a/aluin/sel1_b23/B3 ;
  wire  \t/a/aluin/sel1_b23/B9 ;
  wire  \t/a/aluin/sel1_b24/B2 ;
  wire  \t/a/aluin/sel1_b24/B3 ;
  wire  \t/a/aluin/sel1_b24/B9 ;
  wire  \t/a/aluin/sel1_b25/B2 ;
  wire  \t/a/aluin/sel1_b25/B3 ;
  wire  \t/a/aluin/sel1_b25/B9 ;
  wire  \t/a/aluin/sel1_b26/B2 ;
  wire  \t/a/aluin/sel1_b26/B3 ;
  wire  \t/a/aluin/sel1_b26/B9 ;
  wire  \t/a/aluin/sel1_b27/B2 ;
  wire  \t/a/aluin/sel1_b27/B3 ;
  wire  \t/a/aluin/sel1_b27/B9 ;
  wire  \t/a/aluin/sel1_b28/B2 ;
  wire  \t/a/aluin/sel1_b28/B3 ;
  wire  \t/a/aluin/sel1_b28/B9 ;
  wire  \t/a/aluin/sel1_b29/B2 ;
  wire  \t/a/aluin/sel1_b29/B3 ;
  wire  \t/a/aluin/sel1_b29/B9 ;
  wire  \t/a/aluin/sel1_b3/B6 ;
  wire  \t/a/aluin/sel1_b3/B7 ;
  wire  \t/a/aluin/sel1_b3/B8 ;
  wire  \t/a/aluin/sel1_b3/B9 ;
  wire  \t/a/aluin/sel1_b30/B2 ;
  wire  \t/a/aluin/sel1_b30/B3 ;
  wire  \t/a/aluin/sel1_b30/B9 ;
  wire  \t/a/aluin/sel1_b31/B2 ;
  wire  \t/a/aluin/sel1_b31/B3 ;
  wire  \t/a/aluin/sel1_b31/B9 ;
  wire  \t/a/aluin/sel1_b4/B6 ;
  wire  \t/a/aluin/sel1_b4/B7 ;
  wire  \t/a/aluin/sel1_b4/B8 ;
  wire  \t/a/aluin/sel1_b4/B9 ;
  wire  \t/a/aluin/sel1_b5/B6 ;
  wire  \t/a/aluin/sel1_b5/B7 ;
  wire  \t/a/aluin/sel1_b5/B8 ;
  wire  \t/a/aluin/sel1_b5/B9 ;
  wire  \t/a/aluin/sel1_b6/B6 ;
  wire  \t/a/aluin/sel1_b6/B7 ;
  wire  \t/a/aluin/sel1_b6/B8 ;
  wire  \t/a/aluin/sel1_b6/B9 ;
  wire  \t/a/aluin/sel1_b7/B6 ;
  wire  \t/a/aluin/sel1_b7/B7 ;
  wire  \t/a/aluin/sel1_b7/B8 ;
  wire  \t/a/aluin/sel1_b7/B9 ;
  wire  \t/a/aluin/sel1_b8/B6 ;
  wire  \t/a/aluin/sel1_b8/B7 ;
  wire  \t/a/aluin/sel1_b8/B8 ;
  wire  \t/a/aluin/sel1_b8/B9 ;
  wire  \t/a/aluin/sel1_b9/B6 ;
  wire  \t/a/aluin/sel1_b9/B7 ;
  wire  \t/a/aluin/sel1_b9/B8 ;
  wire  \t/a/aluin/sel1_b9/B9 ;
  wire [31:0] \t/a/condition/JALR_jump_addr ;  // PC.v(257)
  wire [31:0] \t/a/condition/SB_jump_addr ;  // PC.v(260)
  wire [31:0] \t/a/condition/n3 ;
  wire [31:0] \t/a/condition/n5 ;
  wire  \t/a/condition/sel0_b1/B1 ;
  wire  \t/a/condition/sel0_b1/B2 ;
  wire  \t/a/condition/sel0_b10/B1 ;
  wire  \t/a/condition/sel0_b10/B2 ;
  wire  \t/a/condition/sel0_b11/B1 ;
  wire  \t/a/condition/sel0_b11/B2 ;
  wire  \t/a/condition/sel0_b12/B1 ;
  wire  \t/a/condition/sel0_b12/B2 ;
  wire  \t/a/condition/sel0_b13/B2 ;
  wire  \t/a/condition/sel0_b14/B2 ;
  wire  \t/a/condition/sel0_b15/B2 ;
  wire  \t/a/condition/sel0_b16/B2 ;
  wire  \t/a/condition/sel0_b17/B2 ;
  wire  \t/a/condition/sel0_b18/B2 ;
  wire  \t/a/condition/sel0_b19/B2 ;
  wire  \t/a/condition/sel0_b2/B1 ;
  wire  \t/a/condition/sel0_b2/B2 ;
  wire  \t/a/condition/sel0_b20/B2 ;
  wire  \t/a/condition/sel0_b21/B2 ;
  wire  \t/a/condition/sel0_b22/B2 ;
  wire  \t/a/condition/sel0_b23/B2 ;
  wire  \t/a/condition/sel0_b24/B2 ;
  wire  \t/a/condition/sel0_b25/B2 ;
  wire  \t/a/condition/sel0_b26/B2 ;
  wire  \t/a/condition/sel0_b27/B2 ;
  wire  \t/a/condition/sel0_b28/B2 ;
  wire  \t/a/condition/sel0_b29/B2 ;
  wire  \t/a/condition/sel0_b3/B1 ;
  wire  \t/a/condition/sel0_b3/B2 ;
  wire  \t/a/condition/sel0_b30/B2 ;
  wire  \t/a/condition/sel0_b31/B2 ;
  wire  \t/a/condition/sel0_b4/B1 ;
  wire  \t/a/condition/sel0_b4/B2 ;
  wire  \t/a/condition/sel0_b5/B1 ;
  wire  \t/a/condition/sel0_b5/B2 ;
  wire  \t/a/condition/sel0_b6/B1 ;
  wire  \t/a/condition/sel0_b6/B2 ;
  wire  \t/a/condition/sel0_b7/B1 ;
  wire  \t/a/condition/sel0_b7/B2 ;
  wire  \t/a/condition/sel0_b8/B1 ;
  wire  \t/a/condition/sel0_b8/B2 ;
  wire  \t/a/condition/sel0_b9/B1 ;
  wire  \t/a/condition/sel0_b9/B2 ;
  wire  \t/a/condition/sel1/B1 ;
  wire  \t/a/condition/sel1/B2 ;
  wire [6:0] \t/a/if_id/n10 ;
  wire [2:0] \t/a/if_id/n11 ;
  wire [6:0] \t/a/if_id/n12 ;
  wire [4:0] \t/a/if_id/n13 ;
  wire [4:0] \t/a/if_id/n14 ;
  wire [4:0] \t/a/if_id/n15 ;
  wire [31:0] \t/a/instr/n10 ;
  wire [31:0] \t/a/instr/n12 ;
  wire [31:0] \t/a/instr/n14 ;
  wire [31:0] \t/a/instr/n15 ;
  wire [29:0] \t/a/instr/n16 ;
  wire [31:0] \t/a/instr/n17 ;
  wire [31:0] \t/a/instr/n18 ;
  wire [31:0] \t/a/instr/n19 ;
  wire [31:0] \t/a/mem_wb/n5 ;
  wire [31:0] \t/a/memreaddat ;  // cpu.v(67)
  wire [31:0] \t/a/n40 ;
  wire [31:0] \t/a/reg_writedat ;  // cpu.v(68)
  wire [31:0] \t/a/regfile/n46 ;
  wire [31:0] \t/a/regfile/n5 ;
  wire [31:0] \t/a/regfile/n7 ;
  wire [31:0] \t/a/regfile/n8 ;
  wire [31:0] \t/a/regfile/regfile$0$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$1$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$10$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$11$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$12$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$13$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$14$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$15$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$16$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$17$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$18$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$19$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$2$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$20$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$21$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$22$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$23$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$24$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$25$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$26$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$27$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$28$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$29$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$3$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$30$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$31$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$4$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$5$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$6$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$7$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$8$ ;  // register.v(5)
  wire [31:0] \t/a/regfile/regfile$9$ ;  // register.v(5)
  wire [1:0] \t/a/risk_jump/n34 ;
  wire [1:0] \t/a/risk_jump/n49 ;
  wire [1:0] \t/a/risk_jump/rs1_select ;  // PC.v(134)
  wire [1:0] \t/a/risk_jump/rs2_select ;  // PC.v(135)
  wire [31:0] \t/a/unconditional/n2 ;
  wire [31:0] \t/busarbitration/instruction ;  // io.v(35)
  wire [31:0] \t/instruction ;  // top2.v(19)
  wire [31:0] \t/memaddress ;  // top2.v(15)
  wire [31:0] \t/memreaddat ;  // top2.v(16)
  wire [31:0] \t/memstraddress ;  // top2.v(17)
  wire memread;  // __top.v(13)
  wire memwrite_cs;  // __top.v(14)
  wire n0;
  wire n1;
  wire n5;
  wire n6;
  wire n7;
  wire \t/a/ID_LW_block ;  // cpu.v(32)
  wire \t/a/ID_jump_cs ;  // cpu.v(27)
  wire \t/a/ID_jump_risk_block ;  // cpu.v(31)
  wire \t/a/IF_skip_cs ;  // cpu.v(16)
  wire \t/a/WB_regwritecs ;  // cpu.v(69)
  wire \t/a/alu/n0 ;
  wire \t/a/alu/n1 ;
  wire \t/a/alu/n100 ;
  wire \t/a/alu/n101 ;
  wire \t/a/alu/n102 ;
  wire \t/a/alu/n103 ;
  wire \t/a/alu/n104 ;
  wire \t/a/alu/n105 ;
  wire \t/a/alu/n106 ;
  wire \t/a/alu/n107 ;
  wire \t/a/alu/n108 ;
  wire \t/a/alu/n109 ;
  wire \t/a/alu/n110 ;
  wire \t/a/alu/n111 ;
  wire \t/a/alu/n112 ;
  wire \t/a/alu/n113 ;
  wire \t/a/alu/n114 ;
  wire \t/a/alu/n115 ;
  wire \t/a/alu/n116 ;
  wire \t/a/alu/n117 ;
  wire \t/a/alu/n118 ;
  wire \t/a/alu/n119 ;
  wire \t/a/alu/n120 ;
  wire \t/a/alu/n121 ;
  wire \t/a/alu/n122 ;
  wire \t/a/alu/n123 ;
  wire \t/a/alu/n124 ;
  wire \t/a/alu/n125 ;
  wire \t/a/alu/n126 ;
  wire \t/a/alu/n127 ;
  wire \t/a/alu/n128 ;
  wire \t/a/alu/n129 ;
  wire \t/a/alu/n130 ;
  wire \t/a/alu/n131 ;
  wire \t/a/alu/n132 ;
  wire \t/a/alu/n133 ;
  wire \t/a/alu/n134 ;
  wire \t/a/alu/n135 ;
  wire \t/a/alu/n136 ;
  wire \t/a/alu/n137 ;
  wire \t/a/alu/n138 ;
  wire \t/a/alu/n139 ;
  wire \t/a/alu/n140 ;
  wire \t/a/alu/n141 ;
  wire \t/a/alu/n142 ;
  wire \t/a/alu/n143 ;
  wire \t/a/alu/n144 ;
  wire \t/a/alu/n145 ;
  wire \t/a/alu/n146 ;
  wire \t/a/alu/n147 ;
  wire \t/a/alu/n148 ;
  wire \t/a/alu/n149 ;
  wire \t/a/alu/n150 ;
  wire \t/a/alu/n151 ;
  wire \t/a/alu/n152 ;
  wire \t/a/alu/n153 ;
  wire \t/a/alu/n154 ;
  wire \t/a/alu/n155 ;
  wire \t/a/alu/n156 ;
  wire \t/a/alu/n157 ;
  wire \t/a/alu/n158 ;
  wire \t/a/alu/n159 ;
  wire \t/a/alu/n16 ;
  wire \t/a/alu/n160 ;
  wire \t/a/alu/n161 ;
  wire \t/a/alu/n162 ;
  wire \t/a/alu/n163 ;
  wire \t/a/alu/n164 ;
  wire \t/a/alu/n165 ;
  wire \t/a/alu/n166 ;
  wire \t/a/alu/n167 ;
  wire \t/a/alu/n168 ;
  wire \t/a/alu/n169 ;
  wire \t/a/alu/n17 ;
  wire \t/a/alu/n170 ;
  wire \t/a/alu/n171 ;
  wire \t/a/alu/n172 ;
  wire \t/a/alu/n173 ;
  wire \t/a/alu/n174 ;
  wire \t/a/alu/n175 ;
  wire \t/a/alu/n176 ;
  wire \t/a/alu/n177 ;
  wire \t/a/alu/n178 ;
  wire \t/a/alu/n179 ;
  wire \t/a/alu/n18 ;
  wire \t/a/alu/n180 ;
  wire \t/a/alu/n181 ;
  wire \t/a/alu/n182 ;
  wire \t/a/alu/n183 ;
  wire \t/a/alu/n184 ;
  wire \t/a/alu/n185 ;
  wire \t/a/alu/n186 ;
  wire \t/a/alu/n187 ;
  wire \t/a/alu/n188 ;
  wire \t/a/alu/n189 ;
  wire \t/a/alu/n19 ;
  wire \t/a/alu/n190 ;
  wire \t/a/alu/n191 ;
  wire \t/a/alu/n192 ;
  wire \t/a/alu/n193 ;
  wire \t/a/alu/n194 ;
  wire \t/a/alu/n195 ;
  wire \t/a/alu/n196 ;
  wire \t/a/alu/n197 ;
  wire \t/a/alu/n198 ;
  wire \t/a/alu/n199 ;
  wire \t/a/alu/n2 ;
  wire \t/a/alu/n20 ;
  wire \t/a/alu/n200 ;
  wire \t/a/alu/n201 ;
  wire \t/a/alu/n202 ;
  wire \t/a/alu/n203 ;
  wire \t/a/alu/n204 ;
  wire \t/a/alu/n205 ;
  wire \t/a/alu/n206 ;
  wire \t/a/alu/n207 ;
  wire \t/a/alu/n208 ;
  wire \t/a/alu/n209 ;
  wire \t/a/alu/n21 ;
  wire \t/a/alu/n210 ;
  wire \t/a/alu/n211 ;
  wire \t/a/alu/n212 ;
  wire \t/a/alu/n213 ;
  wire \t/a/alu/n214 ;
  wire \t/a/alu/n215 ;
  wire \t/a/alu/n216 ;
  wire \t/a/alu/n217 ;
  wire \t/a/alu/n218 ;
  wire \t/a/alu/n219 ;
  wire \t/a/alu/n22 ;
  wire \t/a/alu/n220 ;
  wire \t/a/alu/n221 ;
  wire \t/a/alu/n222 ;
  wire \t/a/alu/n223 ;
  wire \t/a/alu/n224 ;
  wire \t/a/alu/n225 ;
  wire \t/a/alu/n226 ;
  wire \t/a/alu/n227 ;
  wire \t/a/alu/n228 ;
  wire \t/a/alu/n229 ;
  wire \t/a/alu/n23 ;
  wire \t/a/alu/n230 ;
  wire \t/a/alu/n231 ;
  wire \t/a/alu/n232 ;
  wire \t/a/alu/n233 ;
  wire \t/a/alu/n234 ;
  wire \t/a/alu/n235 ;
  wire \t/a/alu/n236 ;
  wire \t/a/alu/n237 ;
  wire \t/a/alu/n238 ;
  wire \t/a/alu/n239 ;
  wire \t/a/alu/n24 ;
  wire \t/a/alu/n240 ;
  wire \t/a/alu/n241 ;
  wire \t/a/alu/n242 ;
  wire \t/a/alu/n243 ;
  wire \t/a/alu/n244 ;
  wire \t/a/alu/n245 ;
  wire \t/a/alu/n246 ;
  wire \t/a/alu/n247 ;
  wire \t/a/alu/n248 ;
  wire \t/a/alu/n249 ;
  wire \t/a/alu/n25 ;
  wire \t/a/alu/n250 ;
  wire \t/a/alu/n251 ;
  wire \t/a/alu/n252 ;
  wire \t/a/alu/n253 ;
  wire \t/a/alu/n254 ;
  wire \t/a/alu/n255 ;
  wire \t/a/alu/n256 ;
  wire \t/a/alu/n257 ;
  wire \t/a/alu/n258 ;
  wire \t/a/alu/n259 ;
  wire \t/a/alu/n26 ;
  wire \t/a/alu/n260 ;
  wire \t/a/alu/n261 ;
  wire \t/a/alu/n262 ;
  wire \t/a/alu/n263 ;
  wire \t/a/alu/n264 ;
  wire \t/a/alu/n265 ;
  wire \t/a/alu/n266 ;
  wire \t/a/alu/n267 ;
  wire \t/a/alu/n27 ;
  wire \t/a/alu/n28 ;
  wire \t/a/alu/n29 ;
  wire \t/a/alu/n3 ;
  wire \t/a/alu/n30 ;
  wire \t/a/alu/n31 ;
  wire \t/a/alu/n32 ;
  wire \t/a/alu/n33 ;
  wire \t/a/alu/n34 ;
  wire \t/a/alu/n35 ;
  wire \t/a/alu/n36 ;
  wire \t/a/alu/n37 ;
  wire \t/a/alu/n38 ;
  wire \t/a/alu/n39 ;
  wire \t/a/alu/n4 ;
  wire \t/a/alu/n40 ;
  wire \t/a/alu/n41 ;
  wire \t/a/alu/n42 ;
  wire \t/a/alu/n43 ;
  wire \t/a/alu/n44 ;
  wire \t/a/alu/n45 ;
  wire \t/a/alu/n46 ;
  wire \t/a/alu/n47 ;
  wire \t/a/alu/n50 ;
  wire \t/a/alu/n51 ;
  wire \t/a/alu/n52 ;
  wire \t/a/alu/n53 ;
  wire \t/a/alu/n54 ;
  wire \t/a/alu/n55 ;
  wire \t/a/alu/n56 ;
  wire \t/a/alu/n57 ;
  wire \t/a/alu/n58 ;
  wire \t/a/alu/n59 ;
  wire \t/a/alu/n60 ;
  wire \t/a/alu/n61 ;
  wire \t/a/alu/n62 ;
  wire \t/a/alu/n63 ;
  wire \t/a/alu/n64 ;
  wire \t/a/alu/n65 ;
  wire \t/a/alu/n66 ;
  wire \t/a/alu/n67 ;
  wire \t/a/alu/n68 ;
  wire \t/a/alu/n69 ;
  wire \t/a/alu/n70 ;
  wire \t/a/alu/n71 ;
  wire \t/a/alu/n72 ;
  wire \t/a/alu/n73 ;
  wire \t/a/alu/n74 ;
  wire \t/a/alu/n75 ;
  wire \t/a/alu/n76 ;
  wire \t/a/alu/n77 ;
  wire \t/a/alu/n78 ;
  wire \t/a/alu/n79 ;
  wire \t/a/alu/n8 ;
  wire \t/a/alu/n80 ;
  wire \t/a/alu/n81 ;
  wire \t/a/alu/n82 ;
  wire \t/a/alu/n83 ;
  wire \t/a/alu/n84 ;
  wire \t/a/alu/n85 ;
  wire \t/a/alu/n86 ;
  wire \t/a/alu/n87 ;
  wire \t/a/alu/n88 ;
  wire \t/a/alu/n89 ;
  wire \t/a/alu/n9 ;
  wire \t/a/alu/n90 ;
  wire \t/a/alu/n91 ;
  wire \t/a/alu/n92 ;
  wire \t/a/alu/n93 ;
  wire \t/a/alu/n94 ;
  wire \t/a/alu/n95 ;
  wire \t/a/alu/n96 ;
  wire \t/a/alu/n97 ;
  wire \t/a/alu/n98 ;
  wire \t/a/alu/n99 ;
  wire \t/a/aluin/mux3_b1_sel_is_0_o ;
  wire \t/a/aluin/mux3_b1_sel_is_0_o_neg ;
  wire \t/a/aluin/mux4_b1_sel_is_1_o ;
  wire \t/a/aluin/mux4_b1_sel_is_1_o_neg ;
  wire \t/a/aluin/n0 ;
  wire \t/a/aluin/n1 ;
  wire \t/a/aluin/n10 ;
  wire \t/a/aluin/n11 ;
  wire \t/a/aluin/n12 ;
  wire \t/a/aluin/n13 ;
  wire \t/a/aluin/n14 ;
  wire \t/a/aluin/n15 ;
  wire \t/a/aluin/n2 ;
  wire \t/a/aluin/n3 ;
  wire \t/a/aluin/n32 ;
  wire \t/a/aluin/n34 ;
  wire \t/a/aluin/n35 ;
  wire \t/a/aluin/n36 ;
  wire \t/a/aluin/n36_neg ;
  wire \t/a/aluin/n39 ;
  wire \t/a/aluin/n39_neg ;
  wire \t/a/aluin/n4 ;
  wire \t/a/aluin/n5 ;
  wire \t/a/aluin/n6 ;
  wire \t/a/aluin/n7 ;
  wire \t/a/aluin/n8 ;
  wire \t/a/aluin/sel0_b0/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b0/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b1/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b1/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b10/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b10/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b11/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b11/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b12/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b12/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b13/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b13/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b14/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b14/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b15/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b15/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b16/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b16/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b17/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b17/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b18/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b18/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b19/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b19/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b2/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b2/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b20/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b20/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b21/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b21/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b22/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b22/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b23/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b23/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b24/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b24/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b25/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b25/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b26/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b26/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b27/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b27/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b28/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b28/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b29/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b29/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b3/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b3/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b30/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b30/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b31/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b31/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b4/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b4/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b5/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b5/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b6/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b6/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b7/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b7/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b8/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b8/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel0_b9/or_B0_B1_o ;
  wire \t/a/aluin/sel0_b9/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b0/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b0/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b1/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b1/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b10/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b10/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b11/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b11/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b12/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b12/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b12/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b13/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b13/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b13/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b14/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b14/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b14/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b15/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b15/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b15/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b16/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b16/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b16/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b17/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b17/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b17/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b18/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b18/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b18/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b19/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b19/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b19/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b2/or_B5_B6_o ;
  wire \t/a/aluin/sel1_b2/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b2/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b2/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b20/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b20/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b20/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b21/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b21/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b21/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b22/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b22/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b22/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b23/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b23/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b23/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b24/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b24/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b24/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b25/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b25/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b25/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b26/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b26/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b26/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b27/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b27/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b27/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b28/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b28/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b28/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b29/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b29/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b29/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b3/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b3/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b30/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b30/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b30/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b31/or_B2_or_B3_B4_o_o ;
  wire \t/a/aluin/sel1_b31/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b31/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b4/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b4/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b5/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b5/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b6/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b6/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b7/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b7/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b8/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b8/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel1_b9/or_B7_or_B8_B9_o_o ;
  wire \t/a/aluin/sel1_b9/or_B8_B9_o ;
  wire \t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ;
  wire \t/a/aluin/sel2_b0_sel_o ;  // alu.v(89)
  wire \t/a/aluin/sel2_b1_sel_is_1_o ;
  wire \t/a/aluin/sel2_b3_sel_is_3_o ;
  wire \t/a/condition/JALR_jump_cs ;  // PC.v(258)
  wire \t/a/condition/SB_jump_cs ;  // PC.v(261)
  wire \t/a/condition/n0 ;
  wire \t/a/condition/n1 ;
  wire \t/a/condition/n10 ;
  wire \t/a/condition/n11 ;
  wire \t/a/condition/n12 ;
  wire \t/a/condition/n13 ;
  wire \t/a/condition/n7 ;
  wire \t/a/condition/n8 ;
  wire \t/a/condition/n9 ;
  wire \t/a/condition/sel0_b1/or_B1_B2_o ;
  wire \t/a/condition/sel0_b10/or_B1_B2_o ;
  wire \t/a/condition/sel0_b11/or_B1_B2_o ;
  wire \t/a/condition/sel0_b12/or_B1_B2_o ;
  wire \t/a/condition/sel0_b13/or_B1_B2_o ;
  wire \t/a/condition/sel0_b14/or_B1_B2_o ;
  wire \t/a/condition/sel0_b15/or_B1_B2_o ;
  wire \t/a/condition/sel0_b16/or_B1_B2_o ;
  wire \t/a/condition/sel0_b17/or_B1_B2_o ;
  wire \t/a/condition/sel0_b18/or_B1_B2_o ;
  wire \t/a/condition/sel0_b19/or_B1_B2_o ;
  wire \t/a/condition/sel0_b2/or_B1_B2_o ;
  wire \t/a/condition/sel0_b20/or_B1_B2_o ;
  wire \t/a/condition/sel0_b21/or_B1_B2_o ;
  wire \t/a/condition/sel0_b22/or_B1_B2_o ;
  wire \t/a/condition/sel0_b23/or_B1_B2_o ;
  wire \t/a/condition/sel0_b24/or_B1_B2_o ;
  wire \t/a/condition/sel0_b25/or_B1_B2_o ;
  wire \t/a/condition/sel0_b26/or_B1_B2_o ;
  wire \t/a/condition/sel0_b27/or_B1_B2_o ;
  wire \t/a/condition/sel0_b28/or_B1_B2_o ;
  wire \t/a/condition/sel0_b29/or_B1_B2_o ;
  wire \t/a/condition/sel0_b3/or_B1_B2_o ;
  wire \t/a/condition/sel0_b30/or_B1_B2_o ;
  wire \t/a/condition/sel0_b31/or_B1_B2_o ;
  wire \t/a/condition/sel0_b4/or_B1_B2_o ;
  wire \t/a/condition/sel0_b5/or_B1_B2_o ;
  wire \t/a/condition/sel0_b6/or_B1_B2_o ;
  wire \t/a/condition/sel0_b7/or_B1_B2_o ;
  wire \t/a/condition/sel0_b8/or_B1_B2_o ;
  wire \t/a/condition/sel0_b9/or_B1_B2_o ;
  wire \t/a/condition/sel1/or_B1_B2_o ;
  wire \t/a/ex_mem/n0 ;
  wire \t/a/if_id/n1 ;
  wire \t/a/if_id/n2 ;
  wire \t/a/if_id/n3 ;
  wire \t/a/if_id/n4 ;
  wire \t/a/if_id/n5 ;
  wire \t/a/if_id/n6 ;
  wire \t/a/if_id/n7 ;
  wire \t/a/if_id/n9 ;
  wire \t/a/instr/n1 ;
  wire \t/a/instr/n11 ;
  wire \t/a/instr/n1_neg ;
  wire \t/a/instr/n2 ;
  wire \t/a/instr/n20 ;
  wire \t/a/instr/n3 ;
  wire \t/a/instr/n5 ;
  wire \t/a/instr/n7 ;
  wire \t/a/instr/n9 ;
  wire \t/a/mem_wb/n0 ;
  wire \t/a/mem_wb/n1 ;
  wire \t/a/mem_wb/n10 ;
  wire \t/a/mem_wb/n11 ;
  wire \t/a/mem_wb/n12 ;
  wire \t/a/mem_wb/n13 ;
  wire \t/a/mem_wb/n14 ;
  wire \t/a/mem_wb/n2 ;
  wire \t/a/mem_wb/n7 ;
  wire \t/a/mem_wb/n8 ;
  wire \t/a/mem_wb/n9 ;
  wire \t/a/mux3_b0_sel_is_1_o ;
  wire \t/a/mux3_b10_sel_is_3_o ;
  wire \t/a/mux3_b16_sel_is_3_o ;
  wire \t/a/n0 ;
  wire \t/a/n1 ;
  wire \t/a/n10 ;
  wire \t/a/n11 ;
  wire \t/a/n12 ;
  wire \t/a/n13 ;
  wire \t/a/n14 ;
  wire \t/a/n15 ;
  wire \t/a/n16 ;
  wire \t/a/n17 ;
  wire \t/a/n18 ;
  wire \t/a/n19 ;
  wire \t/a/n2 ;
  wire \t/a/n20 ;
  wire \t/a/n21 ;
  wire \t/a/n22 ;
  wire \t/a/n23 ;
  wire \t/a/n24 ;
  wire \t/a/n25 ;
  wire \t/a/n26 ;
  wire \t/a/n27 ;
  wire \t/a/n28 ;
  wire \t/a/n29 ;
  wire \t/a/n3 ;
  wire \t/a/n30 ;
  wire \t/a/n31 ;
  wire \t/a/n32 ;
  wire \t/a/n33 ;
  wire \t/a/n34 ;
  wire \t/a/n35 ;
  wire \t/a/n36 ;
  wire \t/a/n37 ;
  wire \t/a/n4 ;
  wire \t/a/n5 ;
  wire \t/a/n6 ;
  wire \t/a/n7 ;
  wire \t/a/n8 ;
  wire \t/a/n9 ;
  wire \t/a/regfile/mux39_b0_sel_is_3_o ;
  wire \t/a/regfile/mux39_b1000_sel_is_3_o ;
  wire \t/a/regfile/mux39_b100_sel_is_3_o ;
  wire \t/a/regfile/mux39_b128_sel_is_3_o ;
  wire \t/a/regfile/mux39_b160_sel_is_3_o ;
  wire \t/a/regfile/mux39_b192_sel_is_3_o ;
  wire \t/a/regfile/mux39_b224_sel_is_3_o ;
  wire \t/a/regfile/mux39_b256_sel_is_3_o ;
  wire \t/a/regfile/mux39_b288_sel_is_3_o ;
  wire \t/a/regfile/mux39_b320_sel_is_3_o ;
  wire \t/a/regfile/mux39_b32_sel_is_3_o ;
  wire \t/a/regfile/mux39_b352_sel_is_3_o ;
  wire \t/a/regfile/mux39_b384_sel_is_3_o ;
  wire \t/a/regfile/mux39_b416_sel_is_3_o ;
  wire \t/a/regfile/mux39_b448_sel_is_3_o ;
  wire \t/a/regfile/mux39_b480_sel_is_3_o ;
  wire \t/a/regfile/mux39_b512_sel_is_3_o ;
  wire \t/a/regfile/mux39_b544_sel_is_3_o ;
  wire \t/a/regfile/mux39_b576_sel_is_3_o ;
  wire \t/a/regfile/mux39_b608_sel_is_3_o ;
  wire \t/a/regfile/mux39_b640_sel_is_3_o ;
  wire \t/a/regfile/mux39_b64_sel_is_3_o ;
  wire \t/a/regfile/mux39_b672_sel_is_3_o ;
  wire \t/a/regfile/mux39_b704_sel_is_3_o ;
  wire \t/a/regfile/mux39_b736_sel_is_3_o ;
  wire \t/a/regfile/mux39_b768_sel_is_3_o ;
  wire \t/a/regfile/mux39_b800_sel_is_3_o ;
  wire \t/a/regfile/mux39_b832_sel_is_3_o ;
  wire \t/a/regfile/mux39_b864_sel_is_3_o ;
  wire \t/a/regfile/mux39_b896_sel_is_3_o ;
  wire \t/a/regfile/mux39_b928_sel_is_3_o ;
  wire \t/a/regfile/mux39_b960_sel_is_3_o ;
  wire \t/a/regfile/mux4_b0_sel_is_2_o ;
  wire \t/a/regfile/mux4_b0_sel_is_2_o_neg ;
  wire \t/a/regfile/mux5_b0_sel_is_0_o ;
  wire \t/a/regfile/mux6_b0_sel_is_0_o ;
  wire \t/a/regfile/n0 ;
  wire \t/a/regfile/n1 ;
  wire \t/a/regfile/n10 ;
  wire \t/a/regfile/n11 ;
  wire \t/a/regfile/n12 ;
  wire \t/a/regfile/n13 ;
  wire \t/a/regfile/n14 ;
  wire \t/a/regfile/n15 ;
  wire \t/a/regfile/n16 ;
  wire \t/a/regfile/n17 ;
  wire \t/a/regfile/n18 ;
  wire \t/a/regfile/n19 ;
  wire \t/a/regfile/n2 ;
  wire \t/a/regfile/n20 ;
  wire \t/a/regfile/n21 ;
  wire \t/a/regfile/n22 ;
  wire \t/a/regfile/n23 ;
  wire \t/a/regfile/n24 ;
  wire \t/a/regfile/n25 ;
  wire \t/a/regfile/n26 ;
  wire \t/a/regfile/n27 ;
  wire \t/a/regfile/n28 ;
  wire \t/a/regfile/n29 ;
  wire \t/a/regfile/n2_neg ;
  wire \t/a/regfile/n3 ;
  wire \t/a/regfile/n30 ;
  wire \t/a/regfile/n31 ;
  wire \t/a/regfile/n32 ;
  wire \t/a/regfile/n33 ;
  wire \t/a/regfile/n34 ;
  wire \t/a/regfile/n35 ;
  wire \t/a/regfile/n36 ;
  wire \t/a/regfile/n37 ;
  wire \t/a/regfile/n38 ;
  wire \t/a/regfile/n39 ;
  wire \t/a/regfile/n4 ;
  wire \t/a/regfile/n40 ;
  wire \t/a/regfile/n4_neg ;
  wire \t/a/regfile/n6 ;
  wire \t/a/regfile/n80 ;
  wire \t/a/regfile/n9 ;
  wire \t/a/risk_jump/EX_risk ;  // PC.v(137)
  wire \t/a/risk_jump/MEM_risk ;  // PC.v(138)
  wire \t/a/risk_jump/WB_risk ;  // PC.v(139)
  wire \t/a/risk_jump/n1 ;
  wire \t/a/risk_jump/n10 ;
  wire \t/a/risk_jump/n11 ;
  wire \t/a/risk_jump/n12 ;
  wire \t/a/risk_jump/n13 ;
  wire \t/a/risk_jump/n14 ;
  wire \t/a/risk_jump/n15 ;
  wire \t/a/risk_jump/n16 ;
  wire \t/a/risk_jump/n17 ;
  wire \t/a/risk_jump/n19 ;
  wire \t/a/risk_jump/n2 ;
  wire \t/a/risk_jump/n20 ;
  wire \t/a/risk_jump/n21 ;
  wire \t/a/risk_jump/n23 ;
  wire \t/a/risk_jump/n24 ;
  wire \t/a/risk_jump/n25 ;
  wire \t/a/risk_jump/n26 ;
  wire \t/a/risk_jump/n28 ;
  wire \t/a/risk_jump/n29 ;
  wire \t/a/risk_jump/n3 ;
  wire \t/a/risk_jump/n30 ;
  wire \t/a/risk_jump/n31 ;
  wire \t/a/risk_jump/n33 ;
  wire \t/a/risk_jump/n35 ;
  wire \t/a/risk_jump/n36 ;
  wire \t/a/risk_jump/n37 ;
  wire \t/a/risk_jump/n38 ;
  wire \t/a/risk_jump/n39 ;
  wire \t/a/risk_jump/n40 ;
  wire \t/a/risk_jump/n41 ;
  wire \t/a/risk_jump/n42 ;
  wire \t/a/risk_jump/n43 ;
  wire \t/a/risk_jump/n44 ;
  wire \t/a/risk_jump/n45 ;
  wire \t/a/risk_jump/n46 ;
  wire \t/a/risk_jump/n48 ;
  wire \t/a/risk_jump/n5 ;
  wire \t/a/risk_jump/n51 ;
  wire \t/a/risk_jump/n52 ;
  wire \t/a/risk_jump/n53 ;
  wire \t/a/risk_jump/n54 ;
  wire \t/a/risk_jump/n56 ;
  wire \t/a/risk_jump/n57 ;
  wire \t/a/risk_jump/n58 ;
  wire \t/a/risk_jump/n8 ;
  wire \t/a/sel0_b10_sel_o ;  // cpu.v(301)
  wire \t/a/unconditional/mux1_b12_sel_is_0_o ;
  wire \t/a/unconditional/n0 ;
  wire \t/a/unconditional/n0_neg ;
  wire \t/a/unconditional/n1 ;
  wire \t/a/unconditional/n1_neg ;
  wire \t/bus_block ;  // top2.v(13)
  wire \t/busarbitration/mux2_b0_sel_is_2_o ;
  wire \t/busarbitration/mux2_b10_sel_is_2_o ;
  wire \t/busarbitration/mux2_b16_sel_is_2_o ;
  wire \t/busarbitration/mux5_b0_sel_is_3_o ;
  wire \t/busarbitration/mux6_b0_sel_is_3_o ;
  wire \t/busarbitration/mux6_b10_sel_is_3_o ;
  wire \t/busarbitration/mux6_b16_sel_is_3_o ;
  wire \t/busarbitration/n1 ;
  wire \t/busarbitration/n2 ;
  wire \t/busarbitration/n3 ;
  wire \t/instr_read ;  // top2.v(14)
  wire \t/instrnop ;  // top2.v(12)
  wire \t/memread_cs ;  // top2.v(10)

  eq_w1 eq0 (
    .i0(memwrite_cs),
    .i1(1'b1),
    .o(n5));  // __top.v(60)
  eq_w32 eq1 (
    .i0(addr),
    .i1(32'b00000000000000000000010000000010),
    .o(n6));  // __top.v(61)
  reg_ar_as_w1 led_n_reg (
    .clk(clock),
    .d(o_data[0]),
    .en(n7),
    .reset(~rst),
    .set(1'b0),
    .q(led));  // __top.v(63)
  lt_u32_u32 lt0 (
    .ci(1'b0),
    .i0(addr),
    .i1(32'b00000000000000000000000001100000),
    .o(n0));  // __top.v(51)
  EG_LOGIC_DRAM #(
    .ADDR_WIDTH_R(4),
    .ADDR_WIDTH_W(4),
    .DATA_DEPTH_R(12),
    .DATA_DEPTH_W(12),
    .DATA_WIDTH_R(32),
    .DATA_WIDTH_W(32),
    .INIT_FILE("ram.MIF"))
    \m/dram  (
    .di(o_data),
    .raddr(n3),
    .waddr(n2),
    .wclk(clock),
    .we(memwrite_cs),
    .do(i_data));  // ram/ram.v(40)
  binary_mux_s1_w1 mux0_b0 (
    .i0(1'b0),
    .i1(addr[2]),
    .sel(n1),
    .o(n2[0]));  // __top.v(51)
  binary_mux_s1_w1 mux0_b1 (
    .i0(1'b0),
    .i1(addr[3]),
    .sel(n1),
    .o(n2[1]));  // __top.v(51)
  binary_mux_s1_w1 mux0_b2 (
    .i0(1'b0),
    .i1(addr[4]),
    .sel(n1),
    .o(n2[2]));  // __top.v(51)
  binary_mux_s1_w1 mux0_b3 (
    .i0(1'b0),
    .i1(addr[5]),
    .sel(n1),
    .o(n2[3]));  // __top.v(51)
  binary_mux_s1_w1 mux1_b0 (
    .i0(1'b0),
    .i1(addr[2]),
    .sel(memread),
    .o(n3[0]));  // __top.v(55)
  binary_mux_s1_w1 mux1_b1 (
    .i0(1'b0),
    .i1(addr[3]),
    .sel(memread),
    .o(n3[1]));  // __top.v(55)
  binary_mux_s1_w1 mux1_b2 (
    .i0(1'b0),
    .i1(addr[4]),
    .sel(memread),
    .o(n3[2]));  // __top.v(55)
  binary_mux_s1_w1 mux1_b3 (
    .i0(1'b0),
    .i1(addr[5]),
    .sel(memread),
    .o(n3[3]));  // __top.v(55)
  add_pu32_pu32_o32 \t/a/alu/add0  (
    .i0(\t/a/EX_A ),
    .i1({\t/a/EX_B [31:12],\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .o(\t/a/alu/n5 ));  // alu.v(115)
  lt_u32_u32 \t/a/alu/lt0  (
    .ci(1'b0),
    .i0(\t/a/EX_A ),
    .i1({\t/a/EX_B [31:12],\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .o(\t/a/alu/n8 ));  // alu.v(118)
  binary_mux_s4_w1 \t/a/alu/mux0_b0  (
    .i0(\t/a/alu/n5 [0]),
    .i1(\t/a/alu/n7 [0]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [0]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(\t/a/alu/n8 ),
    .i3(\t/a/alu/n8 ),
    .i4(\t/a/alu/n14 [0]),
    .i5(\t/a/alu/n15 [0]),
    .i6(\t/a/alu/n48 [0]),
    .i7(\t/a/alu/n49 [0]),
    .i8(\t/a/alu/n6 [0]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [0]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b1  (
    .i0(\t/a/alu/n5 [1]),
    .i1(\t/a/alu/n7 [1]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [1]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [1]),
    .i5(\t/a/alu/n15 [1]),
    .i6(\t/a/alu/n48 [1]),
    .i7(\t/a/alu/n49 [1]),
    .i8(\t/a/alu/n6 [1]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [1]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b10  (
    .i0(\t/a/alu/n5 [10]),
    .i1(\t/a/alu/n7 [10]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [10]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [10]),
    .i5(\t/a/alu/n15 [10]),
    .i6(\t/a/alu/n48 [10]),
    .i7(\t/a/alu/n49 [10]),
    .i8(\t/a/alu/n6 [10]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [10]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b11  (
    .i0(\t/a/alu/n5 [11]),
    .i1(\t/a/alu/n7 [11]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [11]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [11]),
    .i5(\t/a/alu/n15 [11]),
    .i6(\t/a/alu/n48 [11]),
    .i7(\t/a/alu/n49 [11]),
    .i8(\t/a/alu/n6 [11]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [11]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b12  (
    .i0(\t/a/alu/n5 [12]),
    .i1(\t/a/alu/n7 [12]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [12]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [12]),
    .i5(\t/a/alu/n15 [12]),
    .i6(\t/a/alu/n48 [12]),
    .i7(\t/a/alu/n49 [12]),
    .i8(\t/a/alu/n6 [12]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [12]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b13  (
    .i0(\t/a/alu/n5 [13]),
    .i1(\t/a/alu/n7 [13]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [13]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [13]),
    .i5(\t/a/alu/n15 [13]),
    .i6(\t/a/alu/n48 [13]),
    .i7(\t/a/alu/n49 [13]),
    .i8(\t/a/alu/n6 [13]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [13]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b14  (
    .i0(\t/a/alu/n5 [14]),
    .i1(\t/a/alu/n7 [14]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [14]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [14]),
    .i5(\t/a/alu/n15 [14]),
    .i6(\t/a/alu/n48 [14]),
    .i7(\t/a/alu/n49 [14]),
    .i8(\t/a/alu/n6 [14]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [14]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b15  (
    .i0(\t/a/alu/n5 [15]),
    .i1(\t/a/alu/n7 [15]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [15]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [15]),
    .i5(\t/a/alu/n15 [15]),
    .i6(\t/a/alu/n48 [15]),
    .i7(\t/a/alu/n49 [15]),
    .i8(\t/a/alu/n6 [15]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [15]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b16  (
    .i0(\t/a/alu/n5 [16]),
    .i1(\t/a/alu/n7 [16]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [16]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [16]),
    .i5(\t/a/alu/n15 [16]),
    .i6(\t/a/alu/n48 [16]),
    .i7(\t/a/alu/n49 [16]),
    .i8(\t/a/alu/n6 [16]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [16]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b17  (
    .i0(\t/a/alu/n5 [17]),
    .i1(\t/a/alu/n7 [17]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [17]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [17]),
    .i5(\t/a/alu/n15 [17]),
    .i6(\t/a/alu/n48 [17]),
    .i7(\t/a/alu/n49 [17]),
    .i8(\t/a/alu/n6 [17]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [17]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b18  (
    .i0(\t/a/alu/n5 [18]),
    .i1(\t/a/alu/n7 [18]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [18]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [18]),
    .i5(\t/a/alu/n15 [18]),
    .i6(\t/a/alu/n48 [18]),
    .i7(\t/a/alu/n49 [18]),
    .i8(\t/a/alu/n6 [18]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [18]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b19  (
    .i0(\t/a/alu/n5 [19]),
    .i1(\t/a/alu/n7 [19]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [19]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [19]),
    .i5(\t/a/alu/n15 [19]),
    .i6(\t/a/alu/n48 [19]),
    .i7(\t/a/alu/n49 [19]),
    .i8(\t/a/alu/n6 [19]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [19]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b2  (
    .i0(\t/a/alu/n5 [2]),
    .i1(\t/a/alu/n7 [2]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [2]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [2]),
    .i5(\t/a/alu/n15 [2]),
    .i6(\t/a/alu/n48 [2]),
    .i7(\t/a/alu/n49 [2]),
    .i8(\t/a/alu/n6 [2]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [2]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b20  (
    .i0(\t/a/alu/n5 [20]),
    .i1(\t/a/alu/n7 [20]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [20]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [20]),
    .i5(\t/a/alu/n15 [20]),
    .i6(\t/a/alu/n48 [20]),
    .i7(\t/a/alu/n49 [20]),
    .i8(\t/a/alu/n6 [20]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [20]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b21  (
    .i0(\t/a/alu/n5 [21]),
    .i1(\t/a/alu/n7 [21]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [21]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [21]),
    .i5(\t/a/alu/n15 [21]),
    .i6(\t/a/alu/n48 [21]),
    .i7(\t/a/alu/n49 [21]),
    .i8(\t/a/alu/n6 [21]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [21]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b22  (
    .i0(\t/a/alu/n5 [22]),
    .i1(\t/a/alu/n7 [22]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [22]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [22]),
    .i5(\t/a/alu/n15 [22]),
    .i6(\t/a/alu/n48 [22]),
    .i7(\t/a/alu/n49 [22]),
    .i8(\t/a/alu/n6 [22]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [22]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b23  (
    .i0(\t/a/alu/n5 [23]),
    .i1(\t/a/alu/n7 [23]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [23]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [23]),
    .i5(\t/a/alu/n15 [23]),
    .i6(\t/a/alu/n48 [23]),
    .i7(\t/a/alu/n49 [23]),
    .i8(\t/a/alu/n6 [23]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [23]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b24  (
    .i0(\t/a/alu/n5 [24]),
    .i1(\t/a/alu/n7 [24]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [24]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [24]),
    .i5(\t/a/alu/n15 [24]),
    .i6(\t/a/alu/n48 [24]),
    .i7(\t/a/alu/n49 [24]),
    .i8(\t/a/alu/n6 [24]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [24]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b25  (
    .i0(\t/a/alu/n5 [25]),
    .i1(\t/a/alu/n7 [25]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [25]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [25]),
    .i5(\t/a/alu/n15 [25]),
    .i6(\t/a/alu/n48 [25]),
    .i7(\t/a/alu/n49 [25]),
    .i8(\t/a/alu/n6 [25]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [25]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b26  (
    .i0(\t/a/alu/n5 [26]),
    .i1(\t/a/alu/n7 [26]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [26]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [26]),
    .i5(\t/a/alu/n15 [26]),
    .i6(\t/a/alu/n48 [26]),
    .i7(\t/a/alu/n49 [26]),
    .i8(\t/a/alu/n6 [26]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [26]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b27  (
    .i0(\t/a/alu/n5 [27]),
    .i1(\t/a/alu/n7 [27]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [27]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [27]),
    .i5(\t/a/alu/n15 [27]),
    .i6(\t/a/alu/n48 [27]),
    .i7(\t/a/alu/n49 [27]),
    .i8(\t/a/alu/n6 [27]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [27]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b28  (
    .i0(\t/a/alu/n5 [28]),
    .i1(\t/a/alu/n7 [28]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [28]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [28]),
    .i5(\t/a/alu/n15 [28]),
    .i6(\t/a/alu/n48 [28]),
    .i7(\t/a/alu/n49 [28]),
    .i8(\t/a/alu/n6 [28]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [28]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b29  (
    .i0(\t/a/alu/n5 [29]),
    .i1(\t/a/alu/n7 [29]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [29]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [29]),
    .i5(\t/a/alu/n15 [29]),
    .i6(\t/a/alu/n48 [29]),
    .i7(\t/a/alu/n49 [29]),
    .i8(\t/a/alu/n6 [29]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [29]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b3  (
    .i0(\t/a/alu/n5 [3]),
    .i1(\t/a/alu/n7 [3]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [3]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [3]),
    .i5(\t/a/alu/n15 [3]),
    .i6(\t/a/alu/n48 [3]),
    .i7(\t/a/alu/n49 [3]),
    .i8(\t/a/alu/n6 [3]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [3]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b30  (
    .i0(\t/a/alu/n5 [30]),
    .i1(\t/a/alu/n7 [30]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [30]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [30]),
    .i5(\t/a/alu/n15 [30]),
    .i6(\t/a/alu/n48 [30]),
    .i7(\t/a/alu/n49 [30]),
    .i8(\t/a/alu/n6 [30]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [30]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b31  (
    .i0(\t/a/alu/n5 [31]),
    .i1(\t/a/alu/n7 [31]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [31]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [31]),
    .i5(\t/a/alu/n15 [31]),
    .i6(\t/a/alu/n48 [31]),
    .i7(\t/a/alu/n49 [31]),
    .i8(\t/a/alu/n6 [31]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [31]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b4  (
    .i0(\t/a/alu/n5 [4]),
    .i1(\t/a/alu/n7 [4]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [4]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [4]),
    .i5(\t/a/alu/n15 [4]),
    .i6(\t/a/alu/n48 [4]),
    .i7(\t/a/alu/n49 [4]),
    .i8(\t/a/alu/n6 [4]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [4]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b5  (
    .i0(\t/a/alu/n5 [5]),
    .i1(\t/a/alu/n7 [5]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [5]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [5]),
    .i5(\t/a/alu/n15 [5]),
    .i6(\t/a/alu/n48 [5]),
    .i7(\t/a/alu/n49 [5]),
    .i8(\t/a/alu/n6 [5]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [5]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b6  (
    .i0(\t/a/alu/n5 [6]),
    .i1(\t/a/alu/n7 [6]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [6]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [6]),
    .i5(\t/a/alu/n15 [6]),
    .i6(\t/a/alu/n48 [6]),
    .i7(\t/a/alu/n49 [6]),
    .i8(\t/a/alu/n6 [6]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [6]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b7  (
    .i0(\t/a/alu/n5 [7]),
    .i1(\t/a/alu/n7 [7]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [7]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [7]),
    .i5(\t/a/alu/n15 [7]),
    .i6(\t/a/alu/n48 [7]),
    .i7(\t/a/alu/n49 [7]),
    .i8(\t/a/alu/n6 [7]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [7]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b8  (
    .i0(\t/a/alu/n5 [8]),
    .i1(\t/a/alu/n7 [8]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [8]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [8]),
    .i5(\t/a/alu/n15 [8]),
    .i6(\t/a/alu/n48 [8]),
    .i7(\t/a/alu/n49 [8]),
    .i8(\t/a/alu/n6 [8]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [8]));  // alu.v(126)
  binary_mux_s4_w1 \t/a/alu/mux0_b9  (
    .i0(\t/a/alu/n5 [9]),
    .i1(\t/a/alu/n7 [9]),
    .i10(1'b0),
    .i11(1'b0),
    .i12(1'b0),
    .i13(\t/a/alu/n15 [9]),
    .i14(1'b0),
    .i15(1'b0),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/alu/n14 [9]),
    .i5(\t/a/alu/n15 [9]),
    .i6(\t/a/alu/n48 [9]),
    .i7(\t/a/alu/n49 [9]),
    .i8(\t/a/alu/n6 [9]),
    .i9(1'b0),
    .sel(\t/a/EX_operation ),
    .o(\t/a/aludat [9]));  // alu.v(126)
  add_pu32_mu32_o32 \t/a/alu/sub0  (
    .i0(\t/a/EX_A ),
    .i1({\t/a/EX_B [31:12],\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ,\t/a/EX_B [2],\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ,\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o }),
    .o(\t/a/alu/n6 ));  // alu.v(116)
  AL_MUX \t/a/alu/u1  (
    .i0(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .i1(\t/a/alu/n12 [4]),
    .sel(\t/a/EX_A [4]),
    .o(\t/a/alu/n14 [4]));
  and \t/a/alu/u100  (\t/a/alu/n49 [29], \t/a/EX_A [29], \t/a/EX_B [29]);  // alu.v(124)
  and \t/a/alu/u101  (\t/a/alu/n49 [30], \t/a/EX_A [30], \t/a/EX_B [30]);  // alu.v(124)
  and \t/a/alu/u102  (\t/a/alu/n49 [31], \t/a/EX_A [31], \t/a/EX_B [31]);  // alu.v(124)
  AL_MUX \t/a/alu/u103  (
    .i0(\t/a/EX_A [1]),
    .i1(\t/a/EX_A [2]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n46 ));  // alu.v(121)
  AL_MUX \t/a/alu/u104  (
    .i0(\t/a/EX_A [2]),
    .i1(\t/a/EX_A [3]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n45 ));  // alu.v(121)
  AL_MUX \t/a/alu/u105  (
    .i0(\t/a/EX_A [3]),
    .i1(\t/a/EX_A [4]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n44 ));  // alu.v(121)
  AL_MUX \t/a/alu/u106  (
    .i0(\t/a/EX_A [4]),
    .i1(\t/a/EX_A [5]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n43 ));  // alu.v(121)
  AL_MUX \t/a/alu/u107  (
    .i0(\t/a/EX_A [5]),
    .i1(\t/a/EX_A [6]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n42 ));  // alu.v(121)
  AL_MUX \t/a/alu/u108  (
    .i0(\t/a/EX_A [6]),
    .i1(\t/a/EX_A [7]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n41 ));  // alu.v(121)
  AL_MUX \t/a/alu/u109  (
    .i0(\t/a/EX_A [7]),
    .i1(\t/a/EX_A [8]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n40 ));  // alu.v(121)
  AL_MUX \t/a/alu/u11  (
    .i0(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .i1(\t/a/alu/n12 [0]),
    .sel(\t/a/EX_A [0]),
    .o(\t/a/alu/n14 [0]));
  AL_MUX \t/a/alu/u110  (
    .i0(\t/a/EX_A [8]),
    .i1(\t/a/EX_A [9]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n39 ));  // alu.v(121)
  AL_MUX \t/a/alu/u111  (
    .i0(\t/a/EX_A [9]),
    .i1(\t/a/EX_A [10]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n38 ));  // alu.v(121)
  AL_MUX \t/a/alu/u112  (
    .i0(\t/a/EX_A [10]),
    .i1(\t/a/EX_A [11]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n37 ));  // alu.v(121)
  AL_MUX \t/a/alu/u113  (
    .i0(\t/a/EX_A [11]),
    .i1(\t/a/EX_A [12]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n36 ));  // alu.v(121)
  AL_MUX \t/a/alu/u114  (
    .i0(\t/a/EX_A [12]),
    .i1(\t/a/EX_A [13]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n35 ));  // alu.v(121)
  AL_MUX \t/a/alu/u115  (
    .i0(\t/a/EX_A [13]),
    .i1(\t/a/EX_A [14]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n34 ));  // alu.v(121)
  AL_MUX \t/a/alu/u116  (
    .i0(\t/a/EX_A [14]),
    .i1(\t/a/EX_A [15]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n33 ));  // alu.v(121)
  AL_MUX \t/a/alu/u117  (
    .i0(\t/a/EX_A [15]),
    .i1(\t/a/EX_A [16]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n32 ));  // alu.v(121)
  AL_MUX \t/a/alu/u118  (
    .i0(\t/a/EX_A [16]),
    .i1(\t/a/EX_A [17]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n31 ));  // alu.v(121)
  AL_MUX \t/a/alu/u119  (
    .i0(\t/a/EX_A [17]),
    .i1(\t/a/EX_A [18]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n30 ));  // alu.v(121)
  AL_MUX \t/a/alu/u12  (
    .i0(\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o ),
    .i1(\t/a/alu/n12 [5]),
    .sel(\t/a/EX_A [5]),
    .o(\t/a/alu/n14 [5]));
  AL_MUX \t/a/alu/u120  (
    .i0(\t/a/EX_A [18]),
    .i1(\t/a/EX_A [19]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n29 ));  // alu.v(121)
  AL_MUX \t/a/alu/u121  (
    .i0(\t/a/EX_A [19]),
    .i1(\t/a/EX_A [20]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n28 ));  // alu.v(121)
  AL_MUX \t/a/alu/u122  (
    .i0(\t/a/EX_A [20]),
    .i1(\t/a/EX_A [21]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n27 ));  // alu.v(121)
  AL_MUX \t/a/alu/u123  (
    .i0(\t/a/EX_A [21]),
    .i1(\t/a/EX_A [22]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n26 ));  // alu.v(121)
  AL_MUX \t/a/alu/u124  (
    .i0(\t/a/EX_A [22]),
    .i1(\t/a/EX_A [23]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n25 ));  // alu.v(121)
  AL_MUX \t/a/alu/u125  (
    .i0(\t/a/EX_A [23]),
    .i1(\t/a/EX_A [24]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n24 ));  // alu.v(121)
  AL_MUX \t/a/alu/u126  (
    .i0(\t/a/EX_A [24]),
    .i1(\t/a/EX_A [25]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n23 ));  // alu.v(121)
  AL_MUX \t/a/alu/u127  (
    .i0(\t/a/EX_A [25]),
    .i1(\t/a/EX_A [26]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n22 ));  // alu.v(121)
  AL_MUX \t/a/alu/u128  (
    .i0(\t/a/EX_A [26]),
    .i1(\t/a/EX_A [27]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n21 ));  // alu.v(121)
  AL_MUX \t/a/alu/u129  (
    .i0(\t/a/EX_A [27]),
    .i1(\t/a/EX_A [28]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n20 ));  // alu.v(121)
  AL_MUX \t/a/alu/u13  (
    .i0(\t/a/EX_A [0]),
    .i1(\t/a/EX_A [1]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n47 ));  // alu.v(121)
  AL_MUX \t/a/alu/u130  (
    .i0(\t/a/EX_A [28]),
    .i1(\t/a/EX_A [29]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n19 ));  // alu.v(121)
  AL_MUX \t/a/alu/u131  (
    .i0(\t/a/EX_A [29]),
    .i1(\t/a/EX_A [30]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n18 ));  // alu.v(121)
  AL_MUX \t/a/alu/u132  (
    .i0(\t/a/EX_A [30]),
    .i1(\t/a/EX_A [31]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n17 ));  // alu.v(121)
  AL_MUX \t/a/alu/u133  (
    .i0(\t/a/EX_A [31]),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n16 ));  // alu.v(121)
  AL_MUX \t/a/alu/u134  (
    .i0(\t/a/alu/n47 ),
    .i1(\t/a/alu/n45 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n9 ));  // alu.v(121)
  AL_MUX \t/a/alu/u135  (
    .i0(\t/a/alu/n46 ),
    .i1(\t/a/alu/n44 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n4 ));  // alu.v(121)
  AL_MUX \t/a/alu/u136  (
    .i0(\t/a/alu/n45 ),
    .i1(\t/a/alu/n43 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n2 ));  // alu.v(121)
  AL_MUX \t/a/alu/u137  (
    .i0(\t/a/alu/n44 ),
    .i1(\t/a/alu/n42 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n1 ));  // alu.v(121)
  AL_MUX \t/a/alu/u138  (
    .i0(\t/a/alu/n43 ),
    .i1(\t/a/alu/n41 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n0 ));  // alu.v(121)
  AL_MUX \t/a/alu/u139  (
    .i0(\t/a/alu/n42 ),
    .i1(\t/a/alu/n40 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n3 ));  // alu.v(121)
  and \t/a/alu/u14  (\t/a/alu/n49 [0], \t/a/EX_A [0], \t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o );  // alu.v(124)
  AL_MUX \t/a/alu/u140  (
    .i0(\t/a/alu/n41 ),
    .i1(\t/a/alu/n39 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n81 ));  // alu.v(121)
  AL_MUX \t/a/alu/u141  (
    .i0(\t/a/alu/n40 ),
    .i1(\t/a/alu/n38 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n80 ));  // alu.v(121)
  AL_MUX \t/a/alu/u142  (
    .i0(\t/a/alu/n39 ),
    .i1(\t/a/alu/n37 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n79 ));  // alu.v(121)
  AL_MUX \t/a/alu/u143  (
    .i0(\t/a/alu/n38 ),
    .i1(\t/a/alu/n36 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n78 ));  // alu.v(121)
  AL_MUX \t/a/alu/u144  (
    .i0(\t/a/alu/n37 ),
    .i1(\t/a/alu/n35 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n77 ));  // alu.v(121)
  AL_MUX \t/a/alu/u145  (
    .i0(\t/a/alu/n36 ),
    .i1(\t/a/alu/n34 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n76 ));  // alu.v(121)
  AL_MUX \t/a/alu/u146  (
    .i0(\t/a/alu/n35 ),
    .i1(\t/a/alu/n33 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n75 ));  // alu.v(121)
  AL_MUX \t/a/alu/u147  (
    .i0(\t/a/alu/n34 ),
    .i1(\t/a/alu/n32 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n74 ));  // alu.v(121)
  AL_MUX \t/a/alu/u148  (
    .i0(\t/a/alu/n33 ),
    .i1(\t/a/alu/n31 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n73 ));  // alu.v(121)
  AL_MUX \t/a/alu/u149  (
    .i0(\t/a/alu/n32 ),
    .i1(\t/a/alu/n30 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n72 ));  // alu.v(121)
  AL_MUX \t/a/alu/u15  (
    .i0(\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o ),
    .i1(\t/a/alu/n12 [7]),
    .sel(\t/a/EX_A [7]),
    .o(\t/a/alu/n14 [7]));
  AL_MUX \t/a/alu/u150  (
    .i0(\t/a/alu/n31 ),
    .i1(\t/a/alu/n29 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n71 ));  // alu.v(121)
  AL_MUX \t/a/alu/u151  (
    .i0(\t/a/alu/n30 ),
    .i1(\t/a/alu/n28 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n70 ));  // alu.v(121)
  AL_MUX \t/a/alu/u152  (
    .i0(\t/a/alu/n29 ),
    .i1(\t/a/alu/n27 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n69 ));  // alu.v(121)
  AL_MUX \t/a/alu/u153  (
    .i0(\t/a/alu/n28 ),
    .i1(\t/a/alu/n26 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n68 ));  // alu.v(121)
  AL_MUX \t/a/alu/u154  (
    .i0(\t/a/alu/n27 ),
    .i1(\t/a/alu/n25 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n67 ));  // alu.v(121)
  AL_MUX \t/a/alu/u155  (
    .i0(\t/a/alu/n26 ),
    .i1(\t/a/alu/n24 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n66 ));  // alu.v(121)
  AL_MUX \t/a/alu/u156  (
    .i0(\t/a/alu/n25 ),
    .i1(\t/a/alu/n23 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n65 ));  // alu.v(121)
  AL_MUX \t/a/alu/u157  (
    .i0(\t/a/alu/n24 ),
    .i1(\t/a/alu/n22 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n64 ));  // alu.v(121)
  AL_MUX \t/a/alu/u158  (
    .i0(\t/a/alu/n23 ),
    .i1(\t/a/alu/n21 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n63 ));  // alu.v(121)
  AL_MUX \t/a/alu/u159  (
    .i0(\t/a/alu/n22 ),
    .i1(\t/a/alu/n20 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n62 ));  // alu.v(121)
  AL_MUX \t/a/alu/u16  (
    .i0(\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o ),
    .i1(\t/a/alu/n12 [8]),
    .sel(\t/a/EX_A [8]),
    .o(\t/a/alu/n14 [8]));
  AL_MUX \t/a/alu/u160  (
    .i0(\t/a/alu/n21 ),
    .i1(\t/a/alu/n19 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n61 ));  // alu.v(121)
  AL_MUX \t/a/alu/u161  (
    .i0(\t/a/alu/n20 ),
    .i1(\t/a/alu/n18 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n60 ));  // alu.v(121)
  AL_MUX \t/a/alu/u162  (
    .i0(\t/a/alu/n19 ),
    .i1(\t/a/alu/n17 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n59 ));  // alu.v(121)
  AL_MUX \t/a/alu/u163  (
    .i0(\t/a/alu/n18 ),
    .i1(\t/a/alu/n16 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n58 ));  // alu.v(121)
  AL_MUX \t/a/alu/u164  (
    .i0(\t/a/alu/n17 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n57 ));  // alu.v(121)
  AL_MUX \t/a/alu/u165  (
    .i0(\t/a/alu/n16 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n56 ));  // alu.v(121)
  AL_MUX \t/a/alu/u166  (
    .i0(\t/a/alu/n9 ),
    .i1(\t/a/alu/n0 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n55 ));  // alu.v(121)
  AL_MUX \t/a/alu/u167  (
    .i0(\t/a/alu/n4 ),
    .i1(\t/a/alu/n3 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n54 ));  // alu.v(121)
  AL_MUX \t/a/alu/u168  (
    .i0(\t/a/alu/n2 ),
    .i1(\t/a/alu/n81 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n53 ));  // alu.v(121)
  AL_MUX \t/a/alu/u169  (
    .i0(\t/a/alu/n1 ),
    .i1(\t/a/alu/n80 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n52 ));  // alu.v(121)
  AL_MUX \t/a/alu/u17  (
    .i0(\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o ),
    .i1(\t/a/alu/n12 [9]),
    .sel(\t/a/EX_A [9]),
    .o(\t/a/alu/n14 [9]));
  AL_MUX \t/a/alu/u170  (
    .i0(\t/a/alu/n0 ),
    .i1(\t/a/alu/n79 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n51 ));  // alu.v(121)
  AL_MUX \t/a/alu/u171  (
    .i0(\t/a/alu/n3 ),
    .i1(\t/a/alu/n78 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n50 ));  // alu.v(121)
  AL_MUX \t/a/alu/u172  (
    .i0(\t/a/alu/n81 ),
    .i1(\t/a/alu/n77 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n82 ));  // alu.v(121)
  AL_MUX \t/a/alu/u173  (
    .i0(\t/a/alu/n80 ),
    .i1(\t/a/alu/n76 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n83 ));  // alu.v(121)
  AL_MUX \t/a/alu/u174  (
    .i0(\t/a/alu/n79 ),
    .i1(\t/a/alu/n75 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n84 ));  // alu.v(121)
  AL_MUX \t/a/alu/u175  (
    .i0(\t/a/alu/n78 ),
    .i1(\t/a/alu/n74 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n85 ));  // alu.v(121)
  AL_MUX \t/a/alu/u176  (
    .i0(\t/a/alu/n77 ),
    .i1(\t/a/alu/n73 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n86 ));  // alu.v(121)
  AL_MUX \t/a/alu/u177  (
    .i0(\t/a/alu/n76 ),
    .i1(\t/a/alu/n72 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n87 ));  // alu.v(121)
  AL_MUX \t/a/alu/u178  (
    .i0(\t/a/alu/n75 ),
    .i1(\t/a/alu/n71 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n88 ));  // alu.v(121)
  AL_MUX \t/a/alu/u179  (
    .i0(\t/a/alu/n74 ),
    .i1(\t/a/alu/n70 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n89 ));  // alu.v(121)
  AL_MUX \t/a/alu/u18  (
    .i0(\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o ),
    .i1(\t/a/alu/n12 [10]),
    .sel(\t/a/EX_A [10]),
    .o(\t/a/alu/n14 [10]));
  AL_MUX \t/a/alu/u180  (
    .i0(\t/a/alu/n73 ),
    .i1(\t/a/alu/n69 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n90 ));  // alu.v(121)
  AL_MUX \t/a/alu/u181  (
    .i0(\t/a/alu/n72 ),
    .i1(\t/a/alu/n68 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n91 ));  // alu.v(121)
  AL_MUX \t/a/alu/u182  (
    .i0(\t/a/alu/n71 ),
    .i1(\t/a/alu/n67 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n92 ));  // alu.v(121)
  AL_MUX \t/a/alu/u183  (
    .i0(\t/a/alu/n70 ),
    .i1(\t/a/alu/n66 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n93 ));  // alu.v(121)
  AL_MUX \t/a/alu/u184  (
    .i0(\t/a/alu/n69 ),
    .i1(\t/a/alu/n65 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n94 ));  // alu.v(121)
  AL_MUX \t/a/alu/u185  (
    .i0(\t/a/alu/n68 ),
    .i1(\t/a/alu/n64 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n95 ));  // alu.v(121)
  AL_MUX \t/a/alu/u186  (
    .i0(\t/a/alu/n67 ),
    .i1(\t/a/alu/n63 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n96 ));  // alu.v(121)
  AL_MUX \t/a/alu/u187  (
    .i0(\t/a/alu/n66 ),
    .i1(\t/a/alu/n62 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n97 ));  // alu.v(121)
  AL_MUX \t/a/alu/u188  (
    .i0(\t/a/alu/n65 ),
    .i1(\t/a/alu/n61 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n98 ));  // alu.v(121)
  AL_MUX \t/a/alu/u189  (
    .i0(\t/a/alu/n64 ),
    .i1(\t/a/alu/n60 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n99 ));  // alu.v(121)
  AL_MUX \t/a/alu/u19  (
    .i0(\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o ),
    .i1(\t/a/alu/n12 [11]),
    .sel(\t/a/EX_A [11]),
    .o(\t/a/alu/n14 [11]));
  AL_MUX \t/a/alu/u190  (
    .i0(\t/a/alu/n63 ),
    .i1(\t/a/alu/n59 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n100 ));  // alu.v(121)
  AL_MUX \t/a/alu/u191  (
    .i0(\t/a/alu/n62 ),
    .i1(\t/a/alu/n58 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n101 ));  // alu.v(121)
  AL_MUX \t/a/alu/u192  (
    .i0(\t/a/alu/n61 ),
    .i1(\t/a/alu/n57 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n102 ));  // alu.v(121)
  AL_MUX \t/a/alu/u193  (
    .i0(\t/a/alu/n60 ),
    .i1(\t/a/alu/n56 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n103 ));  // alu.v(121)
  AL_MUX \t/a/alu/u194  (
    .i0(\t/a/alu/n59 ),
    .i1(1'b0),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n104 ));  // alu.v(121)
  AL_MUX \t/a/alu/u195  (
    .i0(\t/a/alu/n58 ),
    .i1(1'b0),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n105 ));  // alu.v(121)
  AL_MUX \t/a/alu/u196  (
    .i0(\t/a/alu/n57 ),
    .i1(1'b0),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n106 ));  // alu.v(121)
  AL_MUX \t/a/alu/u197  (
    .i0(\t/a/alu/n56 ),
    .i1(1'b0),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n107 ));  // alu.v(121)
  AL_MUX \t/a/alu/u198  (
    .i0(\t/a/alu/n55 ),
    .i1(\t/a/alu/n84 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n108 ));  // alu.v(121)
  AL_MUX \t/a/alu/u199  (
    .i0(\t/a/alu/n54 ),
    .i1(\t/a/alu/n85 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n109 ));  // alu.v(121)
  AL_MUX \t/a/alu/u2  (
    .i0(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .i1(\t/a/alu/n12 [3]),
    .sel(\t/a/EX_A [3]),
    .o(\t/a/alu/n14 [3]));
  AL_MUX \t/a/alu/u20  (
    .i0(\t/a/EX_B [12]),
    .i1(\t/a/alu/n12 [12]),
    .sel(\t/a/EX_A [12]),
    .o(\t/a/alu/n14 [12]));
  AL_MUX \t/a/alu/u200  (
    .i0(\t/a/alu/n53 ),
    .i1(\t/a/alu/n86 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n110 ));  // alu.v(121)
  AL_MUX \t/a/alu/u201  (
    .i0(\t/a/alu/n52 ),
    .i1(\t/a/alu/n87 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n111 ));  // alu.v(121)
  AL_MUX \t/a/alu/u202  (
    .i0(\t/a/alu/n51 ),
    .i1(\t/a/alu/n88 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n112 ));  // alu.v(121)
  AL_MUX \t/a/alu/u203  (
    .i0(\t/a/alu/n50 ),
    .i1(\t/a/alu/n89 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n113 ));  // alu.v(121)
  AL_MUX \t/a/alu/u204  (
    .i0(\t/a/alu/n82 ),
    .i1(\t/a/alu/n90 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n114 ));  // alu.v(121)
  AL_MUX \t/a/alu/u205  (
    .i0(\t/a/alu/n83 ),
    .i1(\t/a/alu/n91 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n115 ));  // alu.v(121)
  AL_MUX \t/a/alu/u206  (
    .i0(\t/a/alu/n84 ),
    .i1(\t/a/alu/n92 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n116 ));  // alu.v(121)
  AL_MUX \t/a/alu/u207  (
    .i0(\t/a/alu/n85 ),
    .i1(\t/a/alu/n93 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n117 ));  // alu.v(121)
  AL_MUX \t/a/alu/u208  (
    .i0(\t/a/alu/n86 ),
    .i1(\t/a/alu/n94 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n118 ));  // alu.v(121)
  AL_MUX \t/a/alu/u209  (
    .i0(\t/a/alu/n87 ),
    .i1(\t/a/alu/n95 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n119 ));  // alu.v(121)
  AL_MUX \t/a/alu/u21  (
    .i0(\t/a/EX_B [13]),
    .i1(\t/a/alu/n12 [13]),
    .sel(\t/a/EX_A [13]),
    .o(\t/a/alu/n14 [13]));
  AL_MUX \t/a/alu/u210  (
    .i0(\t/a/alu/n88 ),
    .i1(\t/a/alu/n96 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n120 ));  // alu.v(121)
  AL_MUX \t/a/alu/u211  (
    .i0(\t/a/alu/n89 ),
    .i1(\t/a/alu/n97 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n121 ));  // alu.v(121)
  AL_MUX \t/a/alu/u212  (
    .i0(\t/a/alu/n90 ),
    .i1(\t/a/alu/n98 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n122 ));  // alu.v(121)
  AL_MUX \t/a/alu/u213  (
    .i0(\t/a/alu/n91 ),
    .i1(\t/a/alu/n99 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n123 ));  // alu.v(121)
  AL_MUX \t/a/alu/u214  (
    .i0(\t/a/alu/n92 ),
    .i1(\t/a/alu/n100 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n124 ));  // alu.v(121)
  AL_MUX \t/a/alu/u215  (
    .i0(\t/a/alu/n93 ),
    .i1(\t/a/alu/n101 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n125 ));  // alu.v(121)
  AL_MUX \t/a/alu/u216  (
    .i0(\t/a/alu/n94 ),
    .i1(\t/a/alu/n102 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n126 ));  // alu.v(121)
  AL_MUX \t/a/alu/u217  (
    .i0(\t/a/alu/n95 ),
    .i1(\t/a/alu/n103 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n127 ));  // alu.v(121)
  AL_MUX \t/a/alu/u218  (
    .i0(\t/a/alu/n96 ),
    .i1(\t/a/alu/n104 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n128 ));  // alu.v(121)
  AL_MUX \t/a/alu/u219  (
    .i0(\t/a/alu/n97 ),
    .i1(\t/a/alu/n105 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n129 ));  // alu.v(121)
  AL_MUX \t/a/alu/u22  (
    .i0(\t/a/EX_B [14]),
    .i1(\t/a/alu/n12 [14]),
    .sel(\t/a/EX_A [14]),
    .o(\t/a/alu/n14 [14]));
  AL_MUX \t/a/alu/u220  (
    .i0(\t/a/alu/n98 ),
    .i1(\t/a/alu/n106 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n130 ));  // alu.v(121)
  AL_MUX \t/a/alu/u221  (
    .i0(\t/a/alu/n99 ),
    .i1(\t/a/alu/n107 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n131 ));  // alu.v(121)
  AL_MUX \t/a/alu/u222  (
    .i0(\t/a/alu/n100 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n132 ));  // alu.v(121)
  AL_MUX \t/a/alu/u223  (
    .i0(\t/a/alu/n101 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n133 ));  // alu.v(121)
  AL_MUX \t/a/alu/u224  (
    .i0(\t/a/alu/n102 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n134 ));  // alu.v(121)
  AL_MUX \t/a/alu/u225  (
    .i0(\t/a/alu/n103 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n135 ));  // alu.v(121)
  AL_MUX \t/a/alu/u226  (
    .i0(\t/a/alu/n104 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n136 ));  // alu.v(121)
  AL_MUX \t/a/alu/u227  (
    .i0(\t/a/alu/n105 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n137 ));  // alu.v(121)
  AL_MUX \t/a/alu/u228  (
    .i0(\t/a/alu/n106 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n138 ));  // alu.v(121)
  AL_MUX \t/a/alu/u229  (
    .i0(\t/a/alu/n107 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n139 ));  // alu.v(121)
  AL_MUX \t/a/alu/u23  (
    .i0(\t/a/EX_B [15]),
    .i1(\t/a/alu/n12 [15]),
    .sel(\t/a/EX_A [15]),
    .o(\t/a/alu/n14 [15]));
  AL_MUX \t/a/alu/u230  (
    .i0(\t/a/alu/n108 ),
    .i1(\t/a/alu/n124 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [0]));  // alu.v(121)
  AL_MUX \t/a/alu/u231  (
    .i0(\t/a/alu/n109 ),
    .i1(\t/a/alu/n125 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [1]));  // alu.v(121)
  AL_MUX \t/a/alu/u232  (
    .i0(\t/a/alu/n110 ),
    .i1(\t/a/alu/n126 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [2]));  // alu.v(121)
  AL_MUX \t/a/alu/u233  (
    .i0(\t/a/alu/n111 ),
    .i1(\t/a/alu/n127 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [3]));  // alu.v(121)
  AL_MUX \t/a/alu/u234  (
    .i0(\t/a/alu/n112 ),
    .i1(\t/a/alu/n128 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [4]));  // alu.v(121)
  AL_MUX \t/a/alu/u235  (
    .i0(\t/a/alu/n113 ),
    .i1(\t/a/alu/n129 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [5]));  // alu.v(121)
  AL_MUX \t/a/alu/u236  (
    .i0(\t/a/alu/n114 ),
    .i1(\t/a/alu/n130 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [6]));  // alu.v(121)
  AL_MUX \t/a/alu/u237  (
    .i0(\t/a/alu/n115 ),
    .i1(\t/a/alu/n131 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [7]));  // alu.v(121)
  AL_MUX \t/a/alu/u238  (
    .i0(\t/a/alu/n116 ),
    .i1(\t/a/alu/n132 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [8]));  // alu.v(121)
  AL_MUX \t/a/alu/u239  (
    .i0(\t/a/alu/n117 ),
    .i1(\t/a/alu/n133 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [9]));  // alu.v(121)
  AL_MUX \t/a/alu/u24  (
    .i0(\t/a/EX_B [16]),
    .i1(\t/a/alu/n12 [16]),
    .sel(\t/a/EX_A [16]),
    .o(\t/a/alu/n14 [16]));
  AL_MUX \t/a/alu/u240  (
    .i0(\t/a/alu/n118 ),
    .i1(\t/a/alu/n134 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [10]));  // alu.v(121)
  AL_MUX \t/a/alu/u241  (
    .i0(\t/a/alu/n119 ),
    .i1(\t/a/alu/n135 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [11]));  // alu.v(121)
  AL_MUX \t/a/alu/u242  (
    .i0(\t/a/alu/n120 ),
    .i1(\t/a/alu/n136 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [12]));  // alu.v(121)
  AL_MUX \t/a/alu/u243  (
    .i0(\t/a/alu/n121 ),
    .i1(\t/a/alu/n137 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [13]));  // alu.v(121)
  AL_MUX \t/a/alu/u244  (
    .i0(\t/a/alu/n122 ),
    .i1(\t/a/alu/n138 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [14]));  // alu.v(121)
  AL_MUX \t/a/alu/u245  (
    .i0(\t/a/alu/n123 ),
    .i1(\t/a/alu/n139 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [15]));  // alu.v(121)
  AL_MUX \t/a/alu/u246  (
    .i0(\t/a/alu/n124 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [16]));  // alu.v(121)
  AL_MUX \t/a/alu/u247  (
    .i0(\t/a/alu/n125 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [17]));  // alu.v(121)
  AL_MUX \t/a/alu/u248  (
    .i0(\t/a/alu/n126 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [18]));  // alu.v(121)
  AL_MUX \t/a/alu/u249  (
    .i0(\t/a/alu/n127 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [19]));  // alu.v(121)
  AL_MUX \t/a/alu/u25  (
    .i0(\t/a/EX_B [17]),
    .i1(\t/a/alu/n12 [17]),
    .sel(\t/a/EX_A [17]),
    .o(\t/a/alu/n14 [17]));
  AL_MUX \t/a/alu/u250  (
    .i0(\t/a/alu/n128 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [20]));  // alu.v(121)
  AL_MUX \t/a/alu/u251  (
    .i0(\t/a/alu/n129 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [21]));  // alu.v(121)
  AL_MUX \t/a/alu/u252  (
    .i0(\t/a/alu/n130 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [22]));  // alu.v(121)
  AL_MUX \t/a/alu/u253  (
    .i0(\t/a/alu/n131 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [23]));  // alu.v(121)
  AL_MUX \t/a/alu/u254  (
    .i0(\t/a/alu/n132 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [24]));  // alu.v(121)
  AL_MUX \t/a/alu/u255  (
    .i0(\t/a/alu/n133 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [25]));  // alu.v(121)
  AL_MUX \t/a/alu/u256  (
    .i0(\t/a/alu/n134 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [26]));  // alu.v(121)
  AL_MUX \t/a/alu/u257  (
    .i0(\t/a/alu/n135 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [27]));  // alu.v(121)
  AL_MUX \t/a/alu/u258  (
    .i0(\t/a/alu/n136 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [28]));  // alu.v(121)
  AL_MUX \t/a/alu/u259  (
    .i0(\t/a/alu/n137 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [29]));  // alu.v(121)
  AL_MUX \t/a/alu/u26  (
    .i0(\t/a/EX_B [18]),
    .i1(\t/a/alu/n12 [18]),
    .sel(\t/a/EX_A [18]),
    .o(\t/a/alu/n14 [18]));
  AL_MUX \t/a/alu/u260  (
    .i0(\t/a/alu/n138 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [30]));  // alu.v(121)
  AL_MUX \t/a/alu/u261  (
    .i0(\t/a/alu/n139 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n15 [31]));  // alu.v(121)
  AL_MUX \t/a/alu/u27  (
    .i0(\t/a/EX_B [19]),
    .i1(\t/a/alu/n12 [19]),
    .sel(\t/a/EX_A [19]),
    .o(\t/a/alu/n14 [19]));
  AL_MUX \t/a/alu/u28  (
    .i0(\t/a/EX_B [20]),
    .i1(\t/a/alu/n12 [20]),
    .sel(\t/a/EX_A [20]),
    .o(\t/a/alu/n14 [20]));
  AL_MUX \t/a/alu/u29  (
    .i0(\t/a/EX_B [21]),
    .i1(\t/a/alu/n12 [21]),
    .sel(\t/a/EX_A [21]),
    .o(\t/a/alu/n14 [21]));
  not \t/a/alu/u293  (\t/a/alu/n12 [1], \t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o );  // alu.v(120)
  not \t/a/alu/u294  (\t/a/alu/n12 [2], \t/a/EX_B [2]);  // alu.v(120)
  not \t/a/alu/u295  (\t/a/alu/n12 [3], \t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o );  // alu.v(120)
  not \t/a/alu/u296  (\t/a/alu/n12 [4], \t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o );  // alu.v(120)
  not \t/a/alu/u297  (\t/a/alu/n12 [5], \t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o );  // alu.v(120)
  not \t/a/alu/u298  (\t/a/alu/n12 [6], \t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o );  // alu.v(120)
  not \t/a/alu/u299  (\t/a/alu/n12 [7], \t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o );  // alu.v(120)
  AL_MUX \t/a/alu/u3  (
    .i0(\t/a/EX_B [2]),
    .i1(\t/a/alu/n12 [2]),
    .sel(\t/a/EX_A [2]),
    .o(\t/a/alu/n14 [2]));
  AL_MUX \t/a/alu/u30  (
    .i0(\t/a/EX_B [22]),
    .i1(\t/a/alu/n12 [22]),
    .sel(\t/a/EX_A [22]),
    .o(\t/a/alu/n14 [22]));
  not \t/a/alu/u300  (\t/a/alu/n12 [8], \t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o );  // alu.v(120)
  not \t/a/alu/u301  (\t/a/alu/n12 [9], \t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o );  // alu.v(120)
  not \t/a/alu/u302  (\t/a/alu/n12 [10], \t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o );  // alu.v(120)
  not \t/a/alu/u303  (\t/a/alu/n12 [11], \t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o );  // alu.v(120)
  not \t/a/alu/u304  (\t/a/alu/n12 [12], \t/a/EX_B [12]);  // alu.v(120)
  not \t/a/alu/u305  (\t/a/alu/n12 [13], \t/a/EX_B [13]);  // alu.v(120)
  not \t/a/alu/u306  (\t/a/alu/n12 [14], \t/a/EX_B [14]);  // alu.v(120)
  not \t/a/alu/u307  (\t/a/alu/n12 [15], \t/a/EX_B [15]);  // alu.v(120)
  not \t/a/alu/u308  (\t/a/alu/n12 [16], \t/a/EX_B [16]);  // alu.v(120)
  not \t/a/alu/u309  (\t/a/alu/n12 [17], \t/a/EX_B [17]);  // alu.v(120)
  AL_MUX \t/a/alu/u31  (
    .i0(\t/a/EX_B [23]),
    .i1(\t/a/alu/n12 [23]),
    .sel(\t/a/EX_A [23]),
    .o(\t/a/alu/n14 [23]));
  not \t/a/alu/u310  (\t/a/alu/n12 [18], \t/a/EX_B [18]);  // alu.v(120)
  not \t/a/alu/u311  (\t/a/alu/n12 [19], \t/a/EX_B [19]);  // alu.v(120)
  not \t/a/alu/u312  (\t/a/alu/n12 [20], \t/a/EX_B [20]);  // alu.v(120)
  not \t/a/alu/u313  (\t/a/alu/n12 [21], \t/a/EX_B [21]);  // alu.v(120)
  not \t/a/alu/u314  (\t/a/alu/n12 [22], \t/a/EX_B [22]);  // alu.v(120)
  not \t/a/alu/u315  (\t/a/alu/n12 [23], \t/a/EX_B [23]);  // alu.v(120)
  not \t/a/alu/u316  (\t/a/alu/n12 [24], \t/a/EX_B [24]);  // alu.v(120)
  not \t/a/alu/u317  (\t/a/alu/n12 [25], \t/a/EX_B [25]);  // alu.v(120)
  not \t/a/alu/u318  (\t/a/alu/n12 [26], \t/a/EX_B [26]);  // alu.v(120)
  not \t/a/alu/u319  (\t/a/alu/n12 [27], \t/a/EX_B [27]);  // alu.v(120)
  AL_MUX \t/a/alu/u32  (
    .i0(\t/a/EX_B [24]),
    .i1(\t/a/alu/n12 [24]),
    .sel(\t/a/EX_A [24]),
    .o(\t/a/alu/n14 [24]));
  not \t/a/alu/u320  (\t/a/alu/n12 [28], \t/a/EX_B [28]);  // alu.v(120)
  not \t/a/alu/u321  (\t/a/alu/n12 [29], \t/a/EX_B [29]);  // alu.v(120)
  not \t/a/alu/u322  (\t/a/alu/n12 [30], \t/a/EX_B [30]);  // alu.v(120)
  not \t/a/alu/u323  (\t/a/alu/n12 [31], \t/a/EX_B [31]);  // alu.v(120)
  AL_MUX \t/a/alu/u33  (
    .i0(\t/a/EX_B [25]),
    .i1(\t/a/alu/n12 [25]),
    .sel(\t/a/EX_A [25]),
    .o(\t/a/alu/n14 [25]));
  AL_MUX \t/a/alu/u34  (
    .i0(\t/a/EX_B [26]),
    .i1(\t/a/alu/n12 [26]),
    .sel(\t/a/EX_A [26]),
    .o(\t/a/alu/n14 [26]));
  AL_MUX \t/a/alu/u35  (
    .i0(\t/a/EX_B [27]),
    .i1(\t/a/alu/n12 [27]),
    .sel(\t/a/EX_A [27]),
    .o(\t/a/alu/n14 [27]));
  AL_MUX \t/a/alu/u36  (
    .i0(\t/a/EX_B [28]),
    .i1(\t/a/alu/n12 [28]),
    .sel(\t/a/EX_A [28]),
    .o(\t/a/alu/n14 [28]));
  AL_MUX \t/a/alu/u37  (
    .i0(\t/a/EX_B [29]),
    .i1(\t/a/alu/n12 [29]),
    .sel(\t/a/EX_A [29]),
    .o(\t/a/alu/n14 [29]));
  AL_MUX \t/a/alu/u38  (
    .i0(\t/a/EX_B [30]),
    .i1(\t/a/alu/n12 [30]),
    .sel(\t/a/EX_A [30]),
    .o(\t/a/alu/n14 [30]));
  AL_MUX \t/a/alu/u386  (
    .i0(\t/a/EX_A [30]),
    .i1(\t/a/EX_A [29]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n141 ));  // alu.v(117)
  AL_MUX \t/a/alu/u387  (
    .i0(\t/a/EX_A [29]),
    .i1(\t/a/EX_A [28]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n142 ));  // alu.v(117)
  AL_MUX \t/a/alu/u388  (
    .i0(\t/a/EX_A [28]),
    .i1(\t/a/EX_A [27]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n143 ));  // alu.v(117)
  AL_MUX \t/a/alu/u389  (
    .i0(\t/a/EX_A [27]),
    .i1(\t/a/EX_A [26]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n144 ));  // alu.v(117)
  AL_MUX \t/a/alu/u39  (
    .i0(\t/a/EX_B [31]),
    .i1(\t/a/alu/n12 [31]),
    .sel(\t/a/EX_A [31]),
    .o(\t/a/alu/n14 [31]));
  AL_MUX \t/a/alu/u390  (
    .i0(\t/a/EX_A [26]),
    .i1(\t/a/EX_A [25]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n145 ));  // alu.v(117)
  AL_MUX \t/a/alu/u391  (
    .i0(\t/a/EX_A [25]),
    .i1(\t/a/EX_A [24]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n146 ));  // alu.v(117)
  AL_MUX \t/a/alu/u392  (
    .i0(\t/a/EX_A [24]),
    .i1(\t/a/EX_A [23]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n147 ));  // alu.v(117)
  AL_MUX \t/a/alu/u393  (
    .i0(\t/a/EX_A [23]),
    .i1(\t/a/EX_A [22]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n148 ));  // alu.v(117)
  AL_MUX \t/a/alu/u394  (
    .i0(\t/a/EX_A [22]),
    .i1(\t/a/EX_A [21]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n149 ));  // alu.v(117)
  AL_MUX \t/a/alu/u395  (
    .i0(\t/a/EX_A [21]),
    .i1(\t/a/EX_A [20]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n150 ));  // alu.v(117)
  AL_MUX \t/a/alu/u396  (
    .i0(\t/a/EX_A [20]),
    .i1(\t/a/EX_A [19]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n151 ));  // alu.v(117)
  AL_MUX \t/a/alu/u397  (
    .i0(\t/a/EX_A [19]),
    .i1(\t/a/EX_A [18]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n152 ));  // alu.v(117)
  AL_MUX \t/a/alu/u398  (
    .i0(\t/a/EX_A [18]),
    .i1(\t/a/EX_A [17]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n153 ));  // alu.v(117)
  AL_MUX \t/a/alu/u399  (
    .i0(\t/a/EX_A [17]),
    .i1(\t/a/EX_A [16]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n154 ));  // alu.v(117)
  AL_MUX \t/a/alu/u4  (
    .i0(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .i1(\t/a/alu/n12 [1]),
    .sel(\t/a/EX_A [1]),
    .o(\t/a/alu/n14 [1]));
  or \t/a/alu/u40  (\t/a/alu/n48 [0], \t/a/EX_A [0], \t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o );  // alu.v(123)
  AL_MUX \t/a/alu/u400  (
    .i0(\t/a/EX_A [16]),
    .i1(\t/a/EX_A [15]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n155 ));  // alu.v(117)
  AL_MUX \t/a/alu/u401  (
    .i0(\t/a/EX_A [15]),
    .i1(\t/a/EX_A [14]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n156 ));  // alu.v(117)
  AL_MUX \t/a/alu/u402  (
    .i0(\t/a/EX_A [14]),
    .i1(\t/a/EX_A [13]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n157 ));  // alu.v(117)
  AL_MUX \t/a/alu/u403  (
    .i0(\t/a/EX_A [13]),
    .i1(\t/a/EX_A [12]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n158 ));  // alu.v(117)
  AL_MUX \t/a/alu/u404  (
    .i0(\t/a/EX_A [12]),
    .i1(\t/a/EX_A [11]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n159 ));  // alu.v(117)
  AL_MUX \t/a/alu/u405  (
    .i0(\t/a/EX_A [11]),
    .i1(\t/a/EX_A [10]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n160 ));  // alu.v(117)
  AL_MUX \t/a/alu/u406  (
    .i0(\t/a/EX_A [10]),
    .i1(\t/a/EX_A [9]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n161 ));  // alu.v(117)
  AL_MUX \t/a/alu/u407  (
    .i0(\t/a/EX_A [9]),
    .i1(\t/a/EX_A [8]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n162 ));  // alu.v(117)
  AL_MUX \t/a/alu/u408  (
    .i0(\t/a/EX_A [8]),
    .i1(\t/a/EX_A [7]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n163 ));  // alu.v(117)
  AL_MUX \t/a/alu/u409  (
    .i0(\t/a/EX_A [7]),
    .i1(\t/a/EX_A [6]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n164 ));  // alu.v(117)
  or \t/a/alu/u41  (\t/a/alu/n48 [1], \t/a/EX_A [1], \t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o );  // alu.v(123)
  AL_MUX \t/a/alu/u410  (
    .i0(\t/a/EX_A [6]),
    .i1(\t/a/EX_A [5]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n165 ));  // alu.v(117)
  AL_MUX \t/a/alu/u411  (
    .i0(\t/a/EX_A [5]),
    .i1(\t/a/EX_A [4]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n166 ));  // alu.v(117)
  AL_MUX \t/a/alu/u412  (
    .i0(\t/a/EX_A [4]),
    .i1(\t/a/EX_A [3]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n167 ));  // alu.v(117)
  AL_MUX \t/a/alu/u413  (
    .i0(\t/a/EX_A [3]),
    .i1(\t/a/EX_A [2]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n168 ));  // alu.v(117)
  AL_MUX \t/a/alu/u414  (
    .i0(\t/a/EX_A [2]),
    .i1(\t/a/EX_A [1]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n169 ));  // alu.v(117)
  AL_MUX \t/a/alu/u415  (
    .i0(\t/a/EX_A [1]),
    .i1(\t/a/EX_A [0]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n170 ));  // alu.v(117)
  AL_MUX \t/a/alu/u416  (
    .i0(\t/a/EX_A [0]),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n171 ));  // alu.v(117)
  AL_MUX \t/a/alu/u417  (
    .i0(\t/a/alu/n140 ),
    .i1(\t/a/alu/n142 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n172 ));  // alu.v(117)
  AL_MUX \t/a/alu/u418  (
    .i0(\t/a/alu/n141 ),
    .i1(\t/a/alu/n143 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n173 ));  // alu.v(117)
  AL_MUX \t/a/alu/u419  (
    .i0(\t/a/alu/n142 ),
    .i1(\t/a/alu/n144 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n174 ));  // alu.v(117)
  or \t/a/alu/u42  (\t/a/alu/n48 [2], \t/a/EX_A [2], \t/a/EX_B [2]);  // alu.v(123)
  AL_MUX \t/a/alu/u420  (
    .i0(\t/a/alu/n143 ),
    .i1(\t/a/alu/n145 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n175 ));  // alu.v(117)
  AL_MUX \t/a/alu/u421  (
    .i0(\t/a/alu/n144 ),
    .i1(\t/a/alu/n146 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n176 ));  // alu.v(117)
  AL_MUX \t/a/alu/u422  (
    .i0(\t/a/alu/n145 ),
    .i1(\t/a/alu/n147 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n177 ));  // alu.v(117)
  AL_MUX \t/a/alu/u423  (
    .i0(\t/a/alu/n146 ),
    .i1(\t/a/alu/n148 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n178 ));  // alu.v(117)
  AL_MUX \t/a/alu/u424  (
    .i0(\t/a/alu/n147 ),
    .i1(\t/a/alu/n149 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n179 ));  // alu.v(117)
  AL_MUX \t/a/alu/u425  (
    .i0(\t/a/alu/n148 ),
    .i1(\t/a/alu/n150 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n180 ));  // alu.v(117)
  AL_MUX \t/a/alu/u426  (
    .i0(\t/a/alu/n149 ),
    .i1(\t/a/alu/n151 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n181 ));  // alu.v(117)
  AL_MUX \t/a/alu/u427  (
    .i0(\t/a/alu/n150 ),
    .i1(\t/a/alu/n152 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n182 ));  // alu.v(117)
  AL_MUX \t/a/alu/u428  (
    .i0(\t/a/alu/n151 ),
    .i1(\t/a/alu/n153 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n183 ));  // alu.v(117)
  AL_MUX \t/a/alu/u429  (
    .i0(\t/a/alu/n152 ),
    .i1(\t/a/alu/n154 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n184 ));  // alu.v(117)
  or \t/a/alu/u43  (\t/a/alu/n48 [3], \t/a/EX_A [3], \t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o );  // alu.v(123)
  AL_MUX \t/a/alu/u430  (
    .i0(\t/a/alu/n153 ),
    .i1(\t/a/alu/n155 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n185 ));  // alu.v(117)
  AL_MUX \t/a/alu/u431  (
    .i0(\t/a/alu/n154 ),
    .i1(\t/a/alu/n156 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n186 ));  // alu.v(117)
  AL_MUX \t/a/alu/u432  (
    .i0(\t/a/alu/n155 ),
    .i1(\t/a/alu/n157 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n187 ));  // alu.v(117)
  AL_MUX \t/a/alu/u433  (
    .i0(\t/a/alu/n156 ),
    .i1(\t/a/alu/n158 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n188 ));  // alu.v(117)
  AL_MUX \t/a/alu/u434  (
    .i0(\t/a/alu/n157 ),
    .i1(\t/a/alu/n159 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n189 ));  // alu.v(117)
  AL_MUX \t/a/alu/u435  (
    .i0(\t/a/alu/n158 ),
    .i1(\t/a/alu/n160 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n190 ));  // alu.v(117)
  AL_MUX \t/a/alu/u436  (
    .i0(\t/a/alu/n159 ),
    .i1(\t/a/alu/n161 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n191 ));  // alu.v(117)
  AL_MUX \t/a/alu/u437  (
    .i0(\t/a/alu/n160 ),
    .i1(\t/a/alu/n162 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n192 ));  // alu.v(117)
  AL_MUX \t/a/alu/u438  (
    .i0(\t/a/alu/n161 ),
    .i1(\t/a/alu/n163 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n193 ));  // alu.v(117)
  AL_MUX \t/a/alu/u439  (
    .i0(\t/a/alu/n162 ),
    .i1(\t/a/alu/n164 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n194 ));  // alu.v(117)
  or \t/a/alu/u44  (\t/a/alu/n48 [4], \t/a/EX_A [4], \t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o );  // alu.v(123)
  AL_MUX \t/a/alu/u440  (
    .i0(\t/a/alu/n163 ),
    .i1(\t/a/alu/n165 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n195 ));  // alu.v(117)
  AL_MUX \t/a/alu/u441  (
    .i0(\t/a/alu/n164 ),
    .i1(\t/a/alu/n166 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n196 ));  // alu.v(117)
  AL_MUX \t/a/alu/u442  (
    .i0(\t/a/alu/n165 ),
    .i1(\t/a/alu/n167 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n197 ));  // alu.v(117)
  AL_MUX \t/a/alu/u443  (
    .i0(\t/a/alu/n166 ),
    .i1(\t/a/alu/n168 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n198 ));  // alu.v(117)
  AL_MUX \t/a/alu/u444  (
    .i0(\t/a/alu/n167 ),
    .i1(\t/a/alu/n169 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n199 ));  // alu.v(117)
  AL_MUX \t/a/alu/u445  (
    .i0(\t/a/alu/n168 ),
    .i1(\t/a/alu/n170 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n200 ));  // alu.v(117)
  AL_MUX \t/a/alu/u446  (
    .i0(\t/a/alu/n169 ),
    .i1(\t/a/alu/n171 ),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n201 ));  // alu.v(117)
  AL_MUX \t/a/alu/u447  (
    .i0(\t/a/alu/n170 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n202 ));  // alu.v(117)
  AL_MUX \t/a/alu/u448  (
    .i0(\t/a/alu/n171 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n203 ));  // alu.v(117)
  AL_MUX \t/a/alu/u449  (
    .i0(\t/a/alu/n172 ),
    .i1(\t/a/alu/n176 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n204 ));  // alu.v(117)
  or \t/a/alu/u45  (\t/a/alu/n48 [5], \t/a/EX_A [5], \t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o );  // alu.v(123)
  AL_MUX \t/a/alu/u450  (
    .i0(\t/a/alu/n173 ),
    .i1(\t/a/alu/n177 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n205 ));  // alu.v(117)
  AL_MUX \t/a/alu/u451  (
    .i0(\t/a/alu/n174 ),
    .i1(\t/a/alu/n178 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n206 ));  // alu.v(117)
  AL_MUX \t/a/alu/u452  (
    .i0(\t/a/alu/n175 ),
    .i1(\t/a/alu/n179 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n207 ));  // alu.v(117)
  AL_MUX \t/a/alu/u453  (
    .i0(\t/a/alu/n176 ),
    .i1(\t/a/alu/n180 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n208 ));  // alu.v(117)
  AL_MUX \t/a/alu/u454  (
    .i0(\t/a/alu/n177 ),
    .i1(\t/a/alu/n181 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n209 ));  // alu.v(117)
  AL_MUX \t/a/alu/u455  (
    .i0(\t/a/alu/n178 ),
    .i1(\t/a/alu/n182 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n210 ));  // alu.v(117)
  AL_MUX \t/a/alu/u456  (
    .i0(\t/a/alu/n179 ),
    .i1(\t/a/alu/n183 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n211 ));  // alu.v(117)
  AL_MUX \t/a/alu/u457  (
    .i0(\t/a/alu/n180 ),
    .i1(\t/a/alu/n184 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n212 ));  // alu.v(117)
  AL_MUX \t/a/alu/u458  (
    .i0(\t/a/alu/n181 ),
    .i1(\t/a/alu/n185 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n213 ));  // alu.v(117)
  AL_MUX \t/a/alu/u459  (
    .i0(\t/a/alu/n182 ),
    .i1(\t/a/alu/n186 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n214 ));  // alu.v(117)
  or \t/a/alu/u46  (\t/a/alu/n48 [6], \t/a/EX_A [6], \t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o );  // alu.v(123)
  AL_MUX \t/a/alu/u460  (
    .i0(\t/a/alu/n183 ),
    .i1(\t/a/alu/n187 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n215 ));  // alu.v(117)
  AL_MUX \t/a/alu/u461  (
    .i0(\t/a/alu/n184 ),
    .i1(\t/a/alu/n188 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n216 ));  // alu.v(117)
  AL_MUX \t/a/alu/u462  (
    .i0(\t/a/alu/n185 ),
    .i1(\t/a/alu/n189 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n217 ));  // alu.v(117)
  AL_MUX \t/a/alu/u463  (
    .i0(\t/a/alu/n186 ),
    .i1(\t/a/alu/n190 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n218 ));  // alu.v(117)
  AL_MUX \t/a/alu/u464  (
    .i0(\t/a/alu/n187 ),
    .i1(\t/a/alu/n191 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n219 ));  // alu.v(117)
  AL_MUX \t/a/alu/u465  (
    .i0(\t/a/alu/n188 ),
    .i1(\t/a/alu/n192 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n220 ));  // alu.v(117)
  AL_MUX \t/a/alu/u466  (
    .i0(\t/a/alu/n189 ),
    .i1(\t/a/alu/n193 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n221 ));  // alu.v(117)
  AL_MUX \t/a/alu/u467  (
    .i0(\t/a/alu/n190 ),
    .i1(\t/a/alu/n194 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n222 ));  // alu.v(117)
  AL_MUX \t/a/alu/u468  (
    .i0(\t/a/alu/n191 ),
    .i1(\t/a/alu/n195 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n223 ));  // alu.v(117)
  AL_MUX \t/a/alu/u469  (
    .i0(\t/a/alu/n192 ),
    .i1(\t/a/alu/n196 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n224 ));  // alu.v(117)
  or \t/a/alu/u47  (\t/a/alu/n48 [7], \t/a/EX_A [7], \t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o );  // alu.v(123)
  AL_MUX \t/a/alu/u470  (
    .i0(\t/a/alu/n193 ),
    .i1(\t/a/alu/n197 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n225 ));  // alu.v(117)
  AL_MUX \t/a/alu/u471  (
    .i0(\t/a/alu/n194 ),
    .i1(\t/a/alu/n198 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n226 ));  // alu.v(117)
  AL_MUX \t/a/alu/u472  (
    .i0(\t/a/alu/n195 ),
    .i1(\t/a/alu/n199 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n227 ));  // alu.v(117)
  AL_MUX \t/a/alu/u473  (
    .i0(\t/a/alu/n196 ),
    .i1(\t/a/alu/n200 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n228 ));  // alu.v(117)
  AL_MUX \t/a/alu/u474  (
    .i0(\t/a/alu/n197 ),
    .i1(\t/a/alu/n201 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n229 ));  // alu.v(117)
  AL_MUX \t/a/alu/u475  (
    .i0(\t/a/alu/n198 ),
    .i1(\t/a/alu/n202 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n230 ));  // alu.v(117)
  AL_MUX \t/a/alu/u476  (
    .i0(\t/a/alu/n199 ),
    .i1(\t/a/alu/n203 ),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n231 ));  // alu.v(117)
  AL_MUX \t/a/alu/u477  (
    .i0(\t/a/alu/n200 ),
    .i1(1'b0),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n232 ));  // alu.v(117)
  AL_MUX \t/a/alu/u478  (
    .i0(\t/a/alu/n201 ),
    .i1(1'b0),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n233 ));  // alu.v(117)
  AL_MUX \t/a/alu/u479  (
    .i0(\t/a/alu/n202 ),
    .i1(1'b0),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n234 ));  // alu.v(117)
  or \t/a/alu/u48  (\t/a/alu/n48 [8], \t/a/EX_A [8], \t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o );  // alu.v(123)
  AL_MUX \t/a/alu/u480  (
    .i0(\t/a/alu/n203 ),
    .i1(1'b0),
    .sel(\t/a/EX_B [2]),
    .o(\t/a/alu/n235 ));  // alu.v(117)
  AL_MUX \t/a/alu/u481  (
    .i0(\t/a/alu/n204 ),
    .i1(\t/a/alu/n212 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n236 ));  // alu.v(117)
  AL_MUX \t/a/alu/u482  (
    .i0(\t/a/alu/n205 ),
    .i1(\t/a/alu/n213 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n237 ));  // alu.v(117)
  AL_MUX \t/a/alu/u483  (
    .i0(\t/a/alu/n206 ),
    .i1(\t/a/alu/n214 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n238 ));  // alu.v(117)
  AL_MUX \t/a/alu/u484  (
    .i0(\t/a/alu/n207 ),
    .i1(\t/a/alu/n215 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n239 ));  // alu.v(117)
  AL_MUX \t/a/alu/u485  (
    .i0(\t/a/alu/n208 ),
    .i1(\t/a/alu/n216 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n240 ));  // alu.v(117)
  AL_MUX \t/a/alu/u486  (
    .i0(\t/a/alu/n209 ),
    .i1(\t/a/alu/n217 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n241 ));  // alu.v(117)
  AL_MUX \t/a/alu/u487  (
    .i0(\t/a/alu/n210 ),
    .i1(\t/a/alu/n218 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n242 ));  // alu.v(117)
  AL_MUX \t/a/alu/u488  (
    .i0(\t/a/alu/n211 ),
    .i1(\t/a/alu/n219 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n243 ));  // alu.v(117)
  AL_MUX \t/a/alu/u489  (
    .i0(\t/a/alu/n212 ),
    .i1(\t/a/alu/n220 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n244 ));  // alu.v(117)
  or \t/a/alu/u49  (\t/a/alu/n48 [9], \t/a/EX_A [9], \t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o );  // alu.v(123)
  AL_MUX \t/a/alu/u490  (
    .i0(\t/a/alu/n213 ),
    .i1(\t/a/alu/n221 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n245 ));  // alu.v(117)
  AL_MUX \t/a/alu/u491  (
    .i0(\t/a/alu/n214 ),
    .i1(\t/a/alu/n222 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n246 ));  // alu.v(117)
  AL_MUX \t/a/alu/u492  (
    .i0(\t/a/alu/n215 ),
    .i1(\t/a/alu/n223 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n247 ));  // alu.v(117)
  AL_MUX \t/a/alu/u493  (
    .i0(\t/a/alu/n216 ),
    .i1(\t/a/alu/n224 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n248 ));  // alu.v(117)
  AL_MUX \t/a/alu/u494  (
    .i0(\t/a/alu/n217 ),
    .i1(\t/a/alu/n225 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n249 ));  // alu.v(117)
  AL_MUX \t/a/alu/u495  (
    .i0(\t/a/alu/n218 ),
    .i1(\t/a/alu/n226 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n250 ));  // alu.v(117)
  AL_MUX \t/a/alu/u496  (
    .i0(\t/a/alu/n219 ),
    .i1(\t/a/alu/n227 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n251 ));  // alu.v(117)
  AL_MUX \t/a/alu/u497  (
    .i0(\t/a/alu/n220 ),
    .i1(\t/a/alu/n228 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n252 ));  // alu.v(117)
  AL_MUX \t/a/alu/u498  (
    .i0(\t/a/alu/n221 ),
    .i1(\t/a/alu/n229 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n253 ));  // alu.v(117)
  AL_MUX \t/a/alu/u499  (
    .i0(\t/a/alu/n222 ),
    .i1(\t/a/alu/n230 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n254 ));  // alu.v(117)
  AL_MUX \t/a/alu/u5  (
    .i0(\t/a/EX_A [31]),
    .i1(\t/a/EX_A [30]),
    .sel(\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n140 ));  // alu.v(117)
  or \t/a/alu/u50  (\t/a/alu/n48 [10], \t/a/EX_A [10], \t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o );  // alu.v(123)
  AL_MUX \t/a/alu/u500  (
    .i0(\t/a/alu/n223 ),
    .i1(\t/a/alu/n231 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n255 ));  // alu.v(117)
  AL_MUX \t/a/alu/u501  (
    .i0(\t/a/alu/n224 ),
    .i1(\t/a/alu/n232 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n256 ));  // alu.v(117)
  AL_MUX \t/a/alu/u502  (
    .i0(\t/a/alu/n225 ),
    .i1(\t/a/alu/n233 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n257 ));  // alu.v(117)
  AL_MUX \t/a/alu/u503  (
    .i0(\t/a/alu/n226 ),
    .i1(\t/a/alu/n234 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n258 ));  // alu.v(117)
  AL_MUX \t/a/alu/u504  (
    .i0(\t/a/alu/n227 ),
    .i1(\t/a/alu/n235 ),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n259 ));  // alu.v(117)
  AL_MUX \t/a/alu/u505  (
    .i0(\t/a/alu/n228 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n260 ));  // alu.v(117)
  AL_MUX \t/a/alu/u506  (
    .i0(\t/a/alu/n229 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n261 ));  // alu.v(117)
  AL_MUX \t/a/alu/u507  (
    .i0(\t/a/alu/n230 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n262 ));  // alu.v(117)
  AL_MUX \t/a/alu/u508  (
    .i0(\t/a/alu/n231 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n263 ));  // alu.v(117)
  AL_MUX \t/a/alu/u509  (
    .i0(\t/a/alu/n232 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n264 ));  // alu.v(117)
  or \t/a/alu/u51  (\t/a/alu/n48 [11], \t/a/EX_A [11], \t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o );  // alu.v(123)
  AL_MUX \t/a/alu/u510  (
    .i0(\t/a/alu/n233 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n265 ));  // alu.v(117)
  AL_MUX \t/a/alu/u511  (
    .i0(\t/a/alu/n234 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n266 ));  // alu.v(117)
  AL_MUX \t/a/alu/u512  (
    .i0(\t/a/alu/n235 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n267 ));  // alu.v(117)
  AL_MUX \t/a/alu/u513  (
    .i0(\t/a/alu/n236 ),
    .i1(\t/a/alu/n252 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [31]));  // alu.v(117)
  AL_MUX \t/a/alu/u514  (
    .i0(\t/a/alu/n237 ),
    .i1(\t/a/alu/n253 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [30]));  // alu.v(117)
  AL_MUX \t/a/alu/u515  (
    .i0(\t/a/alu/n238 ),
    .i1(\t/a/alu/n254 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [29]));  // alu.v(117)
  AL_MUX \t/a/alu/u516  (
    .i0(\t/a/alu/n239 ),
    .i1(\t/a/alu/n255 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [28]));  // alu.v(117)
  AL_MUX \t/a/alu/u517  (
    .i0(\t/a/alu/n240 ),
    .i1(\t/a/alu/n256 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [27]));  // alu.v(117)
  AL_MUX \t/a/alu/u518  (
    .i0(\t/a/alu/n241 ),
    .i1(\t/a/alu/n257 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [26]));  // alu.v(117)
  AL_MUX \t/a/alu/u519  (
    .i0(\t/a/alu/n242 ),
    .i1(\t/a/alu/n258 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [25]));  // alu.v(117)
  or \t/a/alu/u52  (\t/a/alu/n48 [12], \t/a/EX_A [12], \t/a/EX_B [12]);  // alu.v(123)
  AL_MUX \t/a/alu/u520  (
    .i0(\t/a/alu/n243 ),
    .i1(\t/a/alu/n259 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [24]));  // alu.v(117)
  AL_MUX \t/a/alu/u521  (
    .i0(\t/a/alu/n244 ),
    .i1(\t/a/alu/n260 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [23]));  // alu.v(117)
  AL_MUX \t/a/alu/u522  (
    .i0(\t/a/alu/n245 ),
    .i1(\t/a/alu/n261 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [22]));  // alu.v(117)
  AL_MUX \t/a/alu/u523  (
    .i0(\t/a/alu/n246 ),
    .i1(\t/a/alu/n262 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [21]));  // alu.v(117)
  AL_MUX \t/a/alu/u524  (
    .i0(\t/a/alu/n247 ),
    .i1(\t/a/alu/n263 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [20]));  // alu.v(117)
  AL_MUX \t/a/alu/u525  (
    .i0(\t/a/alu/n248 ),
    .i1(\t/a/alu/n264 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [19]));  // alu.v(117)
  AL_MUX \t/a/alu/u526  (
    .i0(\t/a/alu/n249 ),
    .i1(\t/a/alu/n265 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [18]));  // alu.v(117)
  AL_MUX \t/a/alu/u527  (
    .i0(\t/a/alu/n250 ),
    .i1(\t/a/alu/n266 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [17]));  // alu.v(117)
  AL_MUX \t/a/alu/u528  (
    .i0(\t/a/alu/n251 ),
    .i1(\t/a/alu/n267 ),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [16]));  // alu.v(117)
  AL_MUX \t/a/alu/u529  (
    .i0(\t/a/alu/n252 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [15]));  // alu.v(117)
  or \t/a/alu/u53  (\t/a/alu/n48 [13], \t/a/EX_A [13], \t/a/EX_B [13]);  // alu.v(123)
  AL_MUX \t/a/alu/u530  (
    .i0(\t/a/alu/n253 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [14]));  // alu.v(117)
  AL_MUX \t/a/alu/u531  (
    .i0(\t/a/alu/n254 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [13]));  // alu.v(117)
  AL_MUX \t/a/alu/u532  (
    .i0(\t/a/alu/n255 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [12]));  // alu.v(117)
  AL_MUX \t/a/alu/u533  (
    .i0(\t/a/alu/n256 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [11]));  // alu.v(117)
  AL_MUX \t/a/alu/u534  (
    .i0(\t/a/alu/n257 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [10]));  // alu.v(117)
  AL_MUX \t/a/alu/u535  (
    .i0(\t/a/alu/n258 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [9]));  // alu.v(117)
  AL_MUX \t/a/alu/u536  (
    .i0(\t/a/alu/n259 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [8]));  // alu.v(117)
  AL_MUX \t/a/alu/u537  (
    .i0(\t/a/alu/n260 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [7]));  // alu.v(117)
  AL_MUX \t/a/alu/u538  (
    .i0(\t/a/alu/n261 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [6]));  // alu.v(117)
  AL_MUX \t/a/alu/u539  (
    .i0(\t/a/alu/n262 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [5]));  // alu.v(117)
  or \t/a/alu/u54  (\t/a/alu/n48 [14], \t/a/EX_A [14], \t/a/EX_B [14]);  // alu.v(123)
  AL_MUX \t/a/alu/u540  (
    .i0(\t/a/alu/n263 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [4]));  // alu.v(117)
  AL_MUX \t/a/alu/u541  (
    .i0(\t/a/alu/n264 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [3]));  // alu.v(117)
  AL_MUX \t/a/alu/u542  (
    .i0(\t/a/alu/n265 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [2]));  // alu.v(117)
  AL_MUX \t/a/alu/u543  (
    .i0(\t/a/alu/n266 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [1]));  // alu.v(117)
  AL_MUX \t/a/alu/u544  (
    .i0(\t/a/alu/n267 ),
    .i1(1'b0),
    .sel(\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o ),
    .o(\t/a/alu/n7 [0]));  // alu.v(117)
  or \t/a/alu/u55  (\t/a/alu/n48 [15], \t/a/EX_A [15], \t/a/EX_B [15]);  // alu.v(123)
  or \t/a/alu/u56  (\t/a/alu/n48 [16], \t/a/EX_A [16], \t/a/EX_B [16]);  // alu.v(123)
  or \t/a/alu/u57  (\t/a/alu/n48 [17], \t/a/EX_A [17], \t/a/EX_B [17]);  // alu.v(123)
  or \t/a/alu/u58  (\t/a/alu/n48 [18], \t/a/EX_A [18], \t/a/EX_B [18]);  // alu.v(123)
  or \t/a/alu/u59  (\t/a/alu/n48 [19], \t/a/EX_A [19], \t/a/EX_B [19]);  // alu.v(123)
  or \t/a/alu/u60  (\t/a/alu/n48 [20], \t/a/EX_A [20], \t/a/EX_B [20]);  // alu.v(123)
  or \t/a/alu/u61  (\t/a/alu/n48 [21], \t/a/EX_A [21], \t/a/EX_B [21]);  // alu.v(123)
  or \t/a/alu/u62  (\t/a/alu/n48 [22], \t/a/EX_A [22], \t/a/EX_B [22]);  // alu.v(123)
  or \t/a/alu/u63  (\t/a/alu/n48 [23], \t/a/EX_A [23], \t/a/EX_B [23]);  // alu.v(123)
  or \t/a/alu/u64  (\t/a/alu/n48 [24], \t/a/EX_A [24], \t/a/EX_B [24]);  // alu.v(123)
  or \t/a/alu/u65  (\t/a/alu/n48 [25], \t/a/EX_A [25], \t/a/EX_B [25]);  // alu.v(123)
  or \t/a/alu/u66  (\t/a/alu/n48 [26], \t/a/EX_A [26], \t/a/EX_B [26]);  // alu.v(123)
  or \t/a/alu/u67  (\t/a/alu/n48 [27], \t/a/EX_A [27], \t/a/EX_B [27]);  // alu.v(123)
  or \t/a/alu/u68  (\t/a/alu/n48 [28], \t/a/EX_A [28], \t/a/EX_B [28]);  // alu.v(123)
  or \t/a/alu/u69  (\t/a/alu/n48 [29], \t/a/EX_A [29], \t/a/EX_B [29]);  // alu.v(123)
  or \t/a/alu/u70  (\t/a/alu/n48 [30], \t/a/EX_A [30], \t/a/EX_B [30]);  // alu.v(123)
  or \t/a/alu/u71  (\t/a/alu/n48 [31], \t/a/EX_A [31], \t/a/EX_B [31]);  // alu.v(123)
  and \t/a/alu/u72  (\t/a/alu/n49 [1], \t/a/EX_A [1], \t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o );  // alu.v(124)
  and \t/a/alu/u73  (\t/a/alu/n49 [2], \t/a/EX_A [2], \t/a/EX_B [2]);  // alu.v(124)
  and \t/a/alu/u74  (\t/a/alu/n49 [3], \t/a/EX_A [3], \t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o );  // alu.v(124)
  and \t/a/alu/u75  (\t/a/alu/n49 [4], \t/a/EX_A [4], \t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o );  // alu.v(124)
  and \t/a/alu/u76  (\t/a/alu/n49 [5], \t/a/EX_A [5], \t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o );  // alu.v(124)
  and \t/a/alu/u77  (\t/a/alu/n49 [6], \t/a/EX_A [6], \t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o );  // alu.v(124)
  and \t/a/alu/u78  (\t/a/alu/n49 [7], \t/a/EX_A [7], \t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o );  // alu.v(124)
  and \t/a/alu/u79  (\t/a/alu/n49 [8], \t/a/EX_A [8], \t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o );  // alu.v(124)
  not \t/a/alu/u8  (\t/a/alu/n12 [0], \t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o );  // alu.v(120)
  and \t/a/alu/u80  (\t/a/alu/n49 [9], \t/a/EX_A [9], \t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o );  // alu.v(124)
  and \t/a/alu/u81  (\t/a/alu/n49 [10], \t/a/EX_A [10], \t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o );  // alu.v(124)
  and \t/a/alu/u82  (\t/a/alu/n49 [11], \t/a/EX_A [11], \t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o );  // alu.v(124)
  and \t/a/alu/u83  (\t/a/alu/n49 [12], \t/a/EX_A [12], \t/a/EX_B [12]);  // alu.v(124)
  and \t/a/alu/u84  (\t/a/alu/n49 [13], \t/a/EX_A [13], \t/a/EX_B [13]);  // alu.v(124)
  and \t/a/alu/u85  (\t/a/alu/n49 [14], \t/a/EX_A [14], \t/a/EX_B [14]);  // alu.v(124)
  and \t/a/alu/u86  (\t/a/alu/n49 [15], \t/a/EX_A [15], \t/a/EX_B [15]);  // alu.v(124)
  and \t/a/alu/u87  (\t/a/alu/n49 [16], \t/a/EX_A [16], \t/a/EX_B [16]);  // alu.v(124)
  and \t/a/alu/u88  (\t/a/alu/n49 [17], \t/a/EX_A [17], \t/a/EX_B [17]);  // alu.v(124)
  and \t/a/alu/u89  (\t/a/alu/n49 [18], \t/a/EX_A [18], \t/a/EX_B [18]);  // alu.v(124)
  AL_MUX \t/a/alu/u9  (
    .i0(\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o ),
    .i1(\t/a/alu/n12 [6]),
    .sel(\t/a/EX_A [6]),
    .o(\t/a/alu/n14 [6]));
  and \t/a/alu/u90  (\t/a/alu/n49 [19], \t/a/EX_A [19], \t/a/EX_B [19]);  // alu.v(124)
  and \t/a/alu/u91  (\t/a/alu/n49 [20], \t/a/EX_A [20], \t/a/EX_B [20]);  // alu.v(124)
  and \t/a/alu/u92  (\t/a/alu/n49 [21], \t/a/EX_A [21], \t/a/EX_B [21]);  // alu.v(124)
  and \t/a/alu/u93  (\t/a/alu/n49 [22], \t/a/EX_A [22], \t/a/EX_B [22]);  // alu.v(124)
  and \t/a/alu/u94  (\t/a/alu/n49 [23], \t/a/EX_A [23], \t/a/EX_B [23]);  // alu.v(124)
  and \t/a/alu/u95  (\t/a/alu/n49 [24], \t/a/EX_A [24], \t/a/EX_B [24]);  // alu.v(124)
  and \t/a/alu/u96  (\t/a/alu/n49 [25], \t/a/EX_A [25], \t/a/EX_B [25]);  // alu.v(124)
  and \t/a/alu/u97  (\t/a/alu/n49 [26], \t/a/EX_A [26], \t/a/EX_B [26]);  // alu.v(124)
  and \t/a/alu/u98  (\t/a/alu/n49 [27], \t/a/EX_A [27], \t/a/EX_B [27]);  // alu.v(124)
  and \t/a/alu/u99  (\t/a/alu/n49 [28], \t/a/EX_A [28], \t/a/EX_B [28]);  // alu.v(124)
  eq_w7 \t/a/aluin/eq0  (
    .i0(\t/a/EX_op ),
    .i1(7'b0110111),
    .o(\t/a/aluin/n1 ));  // alu.v(49)
  eq_w7 \t/a/aluin/eq1  (
    .i0(\t/a/EX_op ),
    .i1(7'b1101111),
    .o(\t/a/aluin/n2 ));  // alu.v(50)
  eq_w3 \t/a/aluin/eq11  (
    .i0(\t/a/EX_fun3 ),
    .i1(3'b000),
    .o(\t/a/aluin/n32 ));  // alu.v(94)
  eq_w7 \t/a/aluin/eq12  (
    .i0(\t/a/EX_fun7 ),
    .i1(7'b0100000),
    .o(\t/a/aluin/n35 ));  // alu.v(94)
  eq_w7 \t/a/aluin/eq2  (
    .i0(\t/a/EX_op ),
    .i1(7'b1100111),
    .o(\t/a/aluin/n3 ));  // alu.v(51)
  eq_w7 \t/a/aluin/eq3  (
    .i0(\t/a/EX_op ),
    .i1(7'b0010111),
    .o(\t/a/aluin/n4 ));  // alu.v(52)
  eq_w3 \t/a/aluin/eq4  (
    .i0(\t/a/EX_fun3 ),
    .i1(3'b001),
    .o(\t/a/aluin/n6 ));  // alu.v(64)
  eq_w3 \t/a/aluin/eq5  (
    .i0(\t/a/EX_fun3 ),
    .i1(3'b101),
    .o(\t/a/aluin/n7 ));  // alu.v(64)
  eq_w7 \t/a/aluin/eq6  (
    .i0(\t/a/EX_op ),
    .i1(7'b0110011),
    .o(\t/a/aluin/n10 ));  // alu.v(60)
  eq_w7 \t/a/aluin/eq7  (
    .i0(\t/a/EX_op ),
    .i1(7'b0000011),
    .o(\t/a/aluin/n11 ));  // alu.v(61)
  eq_w7 \t/a/aluin/eq8  (
    .i0(\t/a/EX_op ),
    .i1(7'b0100011),
    .o(\t/a/aluin/n12 ));  // alu.v(62)
  eq_w7 \t/a/aluin/eq9  (
    .i0(\t/a/EX_op ),
    .i1(7'b0010011),
    .o(\t/a/aluin/n13 ));  // alu.v(63)
  binary_mux_s2_w1 \t/a/aluin/mux0_b0  (
    .i0(\t/a/EX_regdat1 [0]),
    .i1(\t/a/MEM_aludat [0]),
    .i2(\t/a/reg_writedat [0]),
    .i3(\t/a/EX_regdat1 [0]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [0]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b1  (
    .i0(\t/a/EX_regdat1 [1]),
    .i1(\t/a/MEM_aludat [1]),
    .i2(\t/a/reg_writedat [1]),
    .i3(\t/a/EX_regdat1 [1]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [1]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b10  (
    .i0(\t/a/EX_regdat1 [10]),
    .i1(\t/a/MEM_aludat [10]),
    .i2(\t/a/reg_writedat [10]),
    .i3(\t/a/EX_regdat1 [10]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [10]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b11  (
    .i0(\t/a/EX_regdat1 [11]),
    .i1(\t/a/MEM_aludat [11]),
    .i2(\t/a/reg_writedat [11]),
    .i3(\t/a/EX_regdat1 [11]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [11]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b12  (
    .i0(\t/a/EX_regdat1 [12]),
    .i1(\t/a/MEM_aludat [12]),
    .i2(\t/a/reg_writedat [12]),
    .i3(\t/a/EX_regdat1 [12]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [12]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b13  (
    .i0(\t/a/EX_regdat1 [13]),
    .i1(\t/a/MEM_aludat [13]),
    .i2(\t/a/reg_writedat [13]),
    .i3(\t/a/EX_regdat1 [13]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [13]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b14  (
    .i0(\t/a/EX_regdat1 [14]),
    .i1(\t/a/MEM_aludat [14]),
    .i2(\t/a/reg_writedat [14]),
    .i3(\t/a/EX_regdat1 [14]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [14]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b15  (
    .i0(\t/a/EX_regdat1 [15]),
    .i1(\t/a/MEM_aludat [15]),
    .i2(\t/a/reg_writedat [15]),
    .i3(\t/a/EX_regdat1 [15]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [15]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b16  (
    .i0(\t/a/EX_regdat1 [16]),
    .i1(\t/a/MEM_aludat [16]),
    .i2(\t/a/reg_writedat [16]),
    .i3(\t/a/EX_regdat1 [16]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [16]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b17  (
    .i0(\t/a/EX_regdat1 [17]),
    .i1(\t/a/MEM_aludat [17]),
    .i2(\t/a/reg_writedat [17]),
    .i3(\t/a/EX_regdat1 [17]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [17]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b18  (
    .i0(\t/a/EX_regdat1 [18]),
    .i1(\t/a/MEM_aludat [18]),
    .i2(\t/a/reg_writedat [18]),
    .i3(\t/a/EX_regdat1 [18]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [18]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b19  (
    .i0(\t/a/EX_regdat1 [19]),
    .i1(\t/a/MEM_aludat [19]),
    .i2(\t/a/reg_writedat [19]),
    .i3(\t/a/EX_regdat1 [19]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [19]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b2  (
    .i0(\t/a/EX_regdat1 [2]),
    .i1(\t/a/MEM_aludat [2]),
    .i2(\t/a/reg_writedat [2]),
    .i3(\t/a/EX_regdat1 [2]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [2]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b20  (
    .i0(\t/a/EX_regdat1 [20]),
    .i1(\t/a/MEM_aludat [20]),
    .i2(\t/a/reg_writedat [20]),
    .i3(\t/a/EX_regdat1 [20]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [20]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b21  (
    .i0(\t/a/EX_regdat1 [21]),
    .i1(\t/a/MEM_aludat [21]),
    .i2(\t/a/reg_writedat [21]),
    .i3(\t/a/EX_regdat1 [21]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [21]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b22  (
    .i0(\t/a/EX_regdat1 [22]),
    .i1(\t/a/MEM_aludat [22]),
    .i2(\t/a/reg_writedat [22]),
    .i3(\t/a/EX_regdat1 [22]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [22]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b23  (
    .i0(\t/a/EX_regdat1 [23]),
    .i1(\t/a/MEM_aludat [23]),
    .i2(\t/a/reg_writedat [23]),
    .i3(\t/a/EX_regdat1 [23]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [23]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b24  (
    .i0(\t/a/EX_regdat1 [24]),
    .i1(\t/a/MEM_aludat [24]),
    .i2(\t/a/reg_writedat [24]),
    .i3(\t/a/EX_regdat1 [24]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [24]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b25  (
    .i0(\t/a/EX_regdat1 [25]),
    .i1(\t/a/MEM_aludat [25]),
    .i2(\t/a/reg_writedat [25]),
    .i3(\t/a/EX_regdat1 [25]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [25]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b26  (
    .i0(\t/a/EX_regdat1 [26]),
    .i1(\t/a/MEM_aludat [26]),
    .i2(\t/a/reg_writedat [26]),
    .i3(\t/a/EX_regdat1 [26]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [26]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b27  (
    .i0(\t/a/EX_regdat1 [27]),
    .i1(\t/a/MEM_aludat [27]),
    .i2(\t/a/reg_writedat [27]),
    .i3(\t/a/EX_regdat1 [27]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [27]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b28  (
    .i0(\t/a/EX_regdat1 [28]),
    .i1(\t/a/MEM_aludat [28]),
    .i2(\t/a/reg_writedat [28]),
    .i3(\t/a/EX_regdat1 [28]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [28]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b29  (
    .i0(\t/a/EX_regdat1 [29]),
    .i1(\t/a/MEM_aludat [29]),
    .i2(\t/a/reg_writedat [29]),
    .i3(\t/a/EX_regdat1 [29]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [29]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b3  (
    .i0(\t/a/EX_regdat1 [3]),
    .i1(\t/a/MEM_aludat [3]),
    .i2(\t/a/reg_writedat [3]),
    .i3(\t/a/EX_regdat1 [3]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [3]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b30  (
    .i0(\t/a/EX_regdat1 [30]),
    .i1(\t/a/MEM_aludat [30]),
    .i2(\t/a/reg_writedat [30]),
    .i3(\t/a/EX_regdat1 [30]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [30]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b31  (
    .i0(\t/a/EX_regdat1 [31]),
    .i1(\t/a/MEM_aludat [31]),
    .i2(\t/a/reg_writedat [31]),
    .i3(\t/a/EX_regdat1 [31]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [31]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b4  (
    .i0(\t/a/EX_regdat1 [4]),
    .i1(\t/a/MEM_aludat [4]),
    .i2(\t/a/reg_writedat [4]),
    .i3(\t/a/EX_regdat1 [4]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [4]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b5  (
    .i0(\t/a/EX_regdat1 [5]),
    .i1(\t/a/MEM_aludat [5]),
    .i2(\t/a/reg_writedat [5]),
    .i3(\t/a/EX_regdat1 [5]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [5]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b6  (
    .i0(\t/a/EX_regdat1 [6]),
    .i1(\t/a/MEM_aludat [6]),
    .i2(\t/a/reg_writedat [6]),
    .i3(\t/a/EX_regdat1 [6]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [6]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b7  (
    .i0(\t/a/EX_regdat1 [7]),
    .i1(\t/a/MEM_aludat [7]),
    .i2(\t/a/reg_writedat [7]),
    .i3(\t/a/EX_regdat1 [7]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [7]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b8  (
    .i0(\t/a/EX_regdat1 [8]),
    .i1(\t/a/MEM_aludat [8]),
    .i2(\t/a/reg_writedat [8]),
    .i3(\t/a/EX_regdat1 [8]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [8]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux0_b9  (
    .i0(\t/a/EX_regdat1 [9]),
    .i1(\t/a/MEM_aludat [9]),
    .i2(\t/a/reg_writedat [9]),
    .i3(\t/a/EX_regdat1 [9]),
    .sel(\t/a/alu_A_select ),
    .o(\t/a/aluin/o_A1 [9]));  // alu.v(34)
  binary_mux_s2_w1 \t/a/aluin/mux1_b0  (
    .i0(\t/a/EX_regdat2 [0]),
    .i1(\t/a/MEM_aludat [0]),
    .i2(\t/a/reg_writedat [0]),
    .i3(\t/a/EX_regdat2 [0]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [0]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b1  (
    .i0(\t/a/EX_regdat2 [1]),
    .i1(\t/a/MEM_aludat [1]),
    .i2(\t/a/reg_writedat [1]),
    .i3(\t/a/EX_regdat2 [1]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [1]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b10  (
    .i0(\t/a/EX_regdat2 [10]),
    .i1(\t/a/MEM_aludat [10]),
    .i2(\t/a/reg_writedat [10]),
    .i3(\t/a/EX_regdat2 [10]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [10]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b11  (
    .i0(\t/a/EX_regdat2 [11]),
    .i1(\t/a/MEM_aludat [11]),
    .i2(\t/a/reg_writedat [11]),
    .i3(\t/a/EX_regdat2 [11]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [11]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b12  (
    .i0(\t/a/EX_regdat2 [12]),
    .i1(\t/a/MEM_aludat [12]),
    .i2(\t/a/reg_writedat [12]),
    .i3(\t/a/EX_regdat2 [12]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [12]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b13  (
    .i0(\t/a/EX_regdat2 [13]),
    .i1(\t/a/MEM_aludat [13]),
    .i2(\t/a/reg_writedat [13]),
    .i3(\t/a/EX_regdat2 [13]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [13]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b14  (
    .i0(\t/a/EX_regdat2 [14]),
    .i1(\t/a/MEM_aludat [14]),
    .i2(\t/a/reg_writedat [14]),
    .i3(\t/a/EX_regdat2 [14]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [14]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b15  (
    .i0(\t/a/EX_regdat2 [15]),
    .i1(\t/a/MEM_aludat [15]),
    .i2(\t/a/reg_writedat [15]),
    .i3(\t/a/EX_regdat2 [15]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [15]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b16  (
    .i0(\t/a/EX_regdat2 [16]),
    .i1(\t/a/MEM_aludat [16]),
    .i2(\t/a/reg_writedat [16]),
    .i3(\t/a/EX_regdat2 [16]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [16]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b17  (
    .i0(\t/a/EX_regdat2 [17]),
    .i1(\t/a/MEM_aludat [17]),
    .i2(\t/a/reg_writedat [17]),
    .i3(\t/a/EX_regdat2 [17]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [17]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b18  (
    .i0(\t/a/EX_regdat2 [18]),
    .i1(\t/a/MEM_aludat [18]),
    .i2(\t/a/reg_writedat [18]),
    .i3(\t/a/EX_regdat2 [18]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [18]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b19  (
    .i0(\t/a/EX_regdat2 [19]),
    .i1(\t/a/MEM_aludat [19]),
    .i2(\t/a/reg_writedat [19]),
    .i3(\t/a/EX_regdat2 [19]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [19]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b2  (
    .i0(\t/a/EX_regdat2 [2]),
    .i1(\t/a/MEM_aludat [2]),
    .i2(\t/a/reg_writedat [2]),
    .i3(\t/a/EX_regdat2 [2]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [2]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b20  (
    .i0(\t/a/EX_regdat2 [20]),
    .i1(\t/a/MEM_aludat [20]),
    .i2(\t/a/reg_writedat [20]),
    .i3(\t/a/EX_regdat2 [20]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [20]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b21  (
    .i0(\t/a/EX_regdat2 [21]),
    .i1(\t/a/MEM_aludat [21]),
    .i2(\t/a/reg_writedat [21]),
    .i3(\t/a/EX_regdat2 [21]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [21]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b22  (
    .i0(\t/a/EX_regdat2 [22]),
    .i1(\t/a/MEM_aludat [22]),
    .i2(\t/a/reg_writedat [22]),
    .i3(\t/a/EX_regdat2 [22]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [22]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b23  (
    .i0(\t/a/EX_regdat2 [23]),
    .i1(\t/a/MEM_aludat [23]),
    .i2(\t/a/reg_writedat [23]),
    .i3(\t/a/EX_regdat2 [23]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [23]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b24  (
    .i0(\t/a/EX_regdat2 [24]),
    .i1(\t/a/MEM_aludat [24]),
    .i2(\t/a/reg_writedat [24]),
    .i3(\t/a/EX_regdat2 [24]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [24]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b25  (
    .i0(\t/a/EX_regdat2 [25]),
    .i1(\t/a/MEM_aludat [25]),
    .i2(\t/a/reg_writedat [25]),
    .i3(\t/a/EX_regdat2 [25]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [25]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b26  (
    .i0(\t/a/EX_regdat2 [26]),
    .i1(\t/a/MEM_aludat [26]),
    .i2(\t/a/reg_writedat [26]),
    .i3(\t/a/EX_regdat2 [26]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [26]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b27  (
    .i0(\t/a/EX_regdat2 [27]),
    .i1(\t/a/MEM_aludat [27]),
    .i2(\t/a/reg_writedat [27]),
    .i3(\t/a/EX_regdat2 [27]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [27]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b28  (
    .i0(\t/a/EX_regdat2 [28]),
    .i1(\t/a/MEM_aludat [28]),
    .i2(\t/a/reg_writedat [28]),
    .i3(\t/a/EX_regdat2 [28]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [28]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b29  (
    .i0(\t/a/EX_regdat2 [29]),
    .i1(\t/a/MEM_aludat [29]),
    .i2(\t/a/reg_writedat [29]),
    .i3(\t/a/EX_regdat2 [29]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [29]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b3  (
    .i0(\t/a/EX_regdat2 [3]),
    .i1(\t/a/MEM_aludat [3]),
    .i2(\t/a/reg_writedat [3]),
    .i3(\t/a/EX_regdat2 [3]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [3]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b30  (
    .i0(\t/a/EX_regdat2 [30]),
    .i1(\t/a/MEM_aludat [30]),
    .i2(\t/a/reg_writedat [30]),
    .i3(\t/a/EX_regdat2 [30]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [30]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b31  (
    .i0(\t/a/EX_regdat2 [31]),
    .i1(\t/a/MEM_aludat [31]),
    .i2(\t/a/reg_writedat [31]),
    .i3(\t/a/EX_regdat2 [31]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [31]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b4  (
    .i0(\t/a/EX_regdat2 [4]),
    .i1(\t/a/MEM_aludat [4]),
    .i2(\t/a/reg_writedat [4]),
    .i3(\t/a/EX_regdat2 [4]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [4]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b5  (
    .i0(\t/a/EX_regdat2 [5]),
    .i1(\t/a/MEM_aludat [5]),
    .i2(\t/a/reg_writedat [5]),
    .i3(\t/a/EX_regdat2 [5]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [5]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b6  (
    .i0(\t/a/EX_regdat2 [6]),
    .i1(\t/a/MEM_aludat [6]),
    .i2(\t/a/reg_writedat [6]),
    .i3(\t/a/EX_regdat2 [6]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [6]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b7  (
    .i0(\t/a/EX_regdat2 [7]),
    .i1(\t/a/MEM_aludat [7]),
    .i2(\t/a/reg_writedat [7]),
    .i3(\t/a/EX_regdat2 [7]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [7]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b8  (
    .i0(\t/a/EX_regdat2 [8]),
    .i1(\t/a/MEM_aludat [8]),
    .i2(\t/a/reg_writedat [8]),
    .i3(\t/a/EX_regdat2 [8]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [8]));  // alu.v(42)
  binary_mux_s2_w1 \t/a/aluin/mux1_b9  (
    .i0(\t/a/EX_regdat2 [9]),
    .i1(\t/a/MEM_aludat [9]),
    .i2(\t/a/reg_writedat [9]),
    .i3(\t/a/EX_regdat2 [9]),
    .sel(\t/a/alu_B_select ),
    .o(\t/a/aluin/o_B1 [9]));  // alu.v(42)
  binary_mux_s1_w1 \t/a/aluin/mux2_b0  (
    .i0(\t/a/EX_fun3 [0]),
    .i1(1'b1),
    .sel(\t/a/aluin/n39 ),
    .o(\t/a/aluin/n40 [0]));  // alu.v(98)
  binary_mux_s1_w1 \t/a/aluin/mux2_b2  (
    .i0(\t/a/EX_fun3 [2]),
    .i1(1'b1),
    .sel(\t/a/aluin/n39 ),
    .o(\t/a/aluin/n40 [2]));  // alu.v(98)
  binary_mux_s1_w1 \t/a/aluin/mux3_b0  (
    .i0(\t/a/aluin/n40 [0]),
    .i1(1'b0),
    .sel(\t/a/aluin/n36 ),
    .o(\t/a/aluin/n41 [0]));  // alu.v(98)
  and \t/a/aluin/mux3_b1_sel_is_0  (\t/a/aluin/mux3_b1_sel_is_0_o , \t/a/aluin/n36_neg , \t/a/aluin/n39_neg );
  not \t/a/aluin/mux3_b1_sel_is_0_o_inv  (\t/a/aluin/mux3_b1_sel_is_0_o_neg , \t/a/aluin/mux3_b1_sel_is_0_o );
  binary_mux_s1_w1 \t/a/aluin/mux3_b2  (
    .i0(\t/a/aluin/n40 [2]),
    .i1(1'b0),
    .sel(\t/a/aluin/n36 ),
    .o(\t/a/aluin/n41 [2]));  // alu.v(98)
  binary_mux_s1_w1 \t/a/aluin/mux4_b0  (
    .i0(\t/a/EX_fun3 [0]),
    .i1(\t/a/aluin/n41 [0]),
    .sel(\t/a/aluin/sel2_b0_sel_o ),
    .o(\t/a/aluin/operation_R [0]));  // alu.v(100)
  and \t/a/aluin/mux4_b1_sel_is_1  (\t/a/aluin/mux4_b1_sel_is_1_o , \t/a/aluin/sel2_b0_sel_o , \t/a/aluin/mux3_b1_sel_is_0_o_neg );
  not \t/a/aluin/mux4_b1_sel_is_1_o_inv  (\t/a/aluin/mux4_b1_sel_is_1_o_neg , \t/a/aluin/mux4_b1_sel_is_1_o );
  binary_mux_s1_w1 \t/a/aluin/mux4_b2  (
    .i0(\t/a/EX_fun3 [2]),
    .i1(\t/a/aluin/n41 [2]),
    .sel(\t/a/aluin/sel2_b0_sel_o ),
    .o(\t/a/aluin/operation_R [2]));  // alu.v(100)
  binary_mux_s1_w1 \t/a/aluin/mux5_b0  (
    .i0(\t/a/EX_fun7 [0]),
    .i1(1'b0),
    .sel(\t/a/aluin/n8 ),
    .o(\t/a/aluin/n9 [0]));  // alu.v(65)
  binary_mux_s1_w1 \t/a/aluin/mux5_b1  (
    .i0(\t/a/EX_fun7 [1]),
    .i1(1'b0),
    .sel(\t/a/aluin/n8 ),
    .o(\t/a/aluin/n9 [1]));  // alu.v(65)
  binary_mux_s1_w1 \t/a/aluin/mux5_b2  (
    .i0(\t/a/EX_fun7 [2]),
    .i1(1'b0),
    .sel(\t/a/aluin/n8 ),
    .o(\t/a/aluin/n9 [2]));  // alu.v(65)
  binary_mux_s1_w1 \t/a/aluin/mux5_b3  (
    .i0(\t/a/EX_fun7 [3]),
    .i1(1'b0),
    .sel(\t/a/aluin/n8 ),
    .o(\t/a/aluin/n9 [3]));  // alu.v(65)
  binary_mux_s1_w1 \t/a/aluin/mux5_b4  (
    .i0(\t/a/EX_fun7 [4]),
    .i1(1'b0),
    .sel(\t/a/aluin/n8 ),
    .o(\t/a/aluin/n9 [4]));  // alu.v(65)
  binary_mux_s1_w1 \t/a/aluin/mux5_b5  (
    .i0(\t/a/EX_fun7 [5]),
    .i1(1'b0),
    .sel(\t/a/aluin/n8 ),
    .o(\t/a/aluin/n9 [5]));  // alu.v(65)
  binary_mux_s1_w1 \t/a/aluin/mux5_b6  (
    .i0(\t/a/EX_fun7 [6]),
    .i1(1'b0),
    .sel(\t/a/aluin/n8 ),
    .o(\t/a/aluin/n9 [6]));  // alu.v(65)
  not \t/a/aluin/n36_inv  (\t/a/aluin/n36_neg , \t/a/aluin/n36 );
  not \t/a/aluin/n39_inv  (\t/a/aluin/n39_neg , \t/a/aluin/n39 );
  and \t/a/aluin/sel0_b0/and_b0_0  (\t/a/aluin/sel0_b0/B0 , \t/a/aluin/o_A1 [0], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b0/and_b0_1  (\t/a/aluin/sel0_b0/B1 , \t/a/EX_memstraddr [0], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b0/and_b0_2  (\t/a/aluin/sel0_b0/B2 , \t/a/EX_memstraddr [0], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b0/and_b0_3  (\t/a/aluin/sel0_b0/B3 , \t/a/EX_memstraddr [0], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b0/or_B0_B1  (\t/a/aluin/sel0_b0/or_B0_B1_o , \t/a/aluin/sel0_b0/B0 , \t/a/aluin/sel0_b0/B1 );
  or \t/a/aluin/sel0_b0/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b0/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b0/B2 , \t/a/aluin/sel0_b0/B3 );
  or \t/a/aluin/sel0_b0/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [0], \t/a/aluin/sel0_b0/or_B0_B1_o , \t/a/aluin/sel0_b0/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b1/and_b0_0  (\t/a/aluin/sel0_b1/B0 , \t/a/aluin/o_A1 [1], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b1/and_b0_1  (\t/a/aluin/sel0_b1/B1 , \t/a/EX_memstraddr [1], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b1/and_b0_2  (\t/a/aluin/sel0_b1/B2 , \t/a/EX_memstraddr [1], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b1/and_b0_3  (\t/a/aluin/sel0_b1/B3 , \t/a/EX_memstraddr [1], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b1/or_B0_B1  (\t/a/aluin/sel0_b1/or_B0_B1_o , \t/a/aluin/sel0_b1/B0 , \t/a/aluin/sel0_b1/B1 );
  or \t/a/aluin/sel0_b1/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b1/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b1/B2 , \t/a/aluin/sel0_b1/B3 );
  or \t/a/aluin/sel0_b1/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [1], \t/a/aluin/sel0_b1/or_B0_B1_o , \t/a/aluin/sel0_b1/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b10/and_b0_0  (\t/a/aluin/sel0_b10/B0 , \t/a/aluin/o_A1 [10], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b10/and_b0_1  (\t/a/aluin/sel0_b10/B1 , \t/a/EX_memstraddr [10], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b10/and_b0_2  (\t/a/aluin/sel0_b10/B2 , \t/a/EX_memstraddr [10], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b10/and_b0_3  (\t/a/aluin/sel0_b10/B3 , \t/a/EX_memstraddr [10], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b10/or_B0_B1  (\t/a/aluin/sel0_b10/or_B0_B1_o , \t/a/aluin/sel0_b10/B0 , \t/a/aluin/sel0_b10/B1 );
  or \t/a/aluin/sel0_b10/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b10/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b10/B2 , \t/a/aluin/sel0_b10/B3 );
  or \t/a/aluin/sel0_b10/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [10], \t/a/aluin/sel0_b10/or_B0_B1_o , \t/a/aluin/sel0_b10/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b11/and_b0_0  (\t/a/aluin/sel0_b11/B0 , \t/a/aluin/o_A1 [11], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b11/and_b0_1  (\t/a/aluin/sel0_b11/B1 , \t/a/EX_memstraddr [11], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b11/and_b0_2  (\t/a/aluin/sel0_b11/B2 , \t/a/EX_memstraddr [11], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b11/and_b0_3  (\t/a/aluin/sel0_b11/B3 , \t/a/EX_memstraddr [11], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b11/or_B0_B1  (\t/a/aluin/sel0_b11/or_B0_B1_o , \t/a/aluin/sel0_b11/B0 , \t/a/aluin/sel0_b11/B1 );
  or \t/a/aluin/sel0_b11/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b11/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b11/B2 , \t/a/aluin/sel0_b11/B3 );
  or \t/a/aluin/sel0_b11/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [11], \t/a/aluin/sel0_b11/or_B0_B1_o , \t/a/aluin/sel0_b11/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b12/and_b0_0  (\t/a/aluin/sel0_b12/B0 , \t/a/aluin/o_A1 [12], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b12/and_b0_1  (\t/a/aluin/sel0_b12/B1 , \t/a/EX_memstraddr [12], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b12/and_b0_2  (\t/a/aluin/sel0_b12/B2 , \t/a/EX_memstraddr [12], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b12/and_b0_3  (\t/a/aluin/sel0_b12/B3 , \t/a/EX_memstraddr [12], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b12/or_B0_B1  (\t/a/aluin/sel0_b12/or_B0_B1_o , \t/a/aluin/sel0_b12/B0 , \t/a/aluin/sel0_b12/B1 );
  or \t/a/aluin/sel0_b12/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b12/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b12/B2 , \t/a/aluin/sel0_b12/B3 );
  or \t/a/aluin/sel0_b12/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [12], \t/a/aluin/sel0_b12/or_B0_B1_o , \t/a/aluin/sel0_b12/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b13/and_b0_0  (\t/a/aluin/sel0_b13/B0 , \t/a/aluin/o_A1 [13], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b13/and_b0_1  (\t/a/aluin/sel0_b13/B1 , \t/a/EX_memstraddr [13], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b13/and_b0_2  (\t/a/aluin/sel0_b13/B2 , \t/a/EX_memstraddr [13], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b13/and_b0_3  (\t/a/aluin/sel0_b13/B3 , \t/a/EX_memstraddr [13], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b13/or_B0_B1  (\t/a/aluin/sel0_b13/or_B0_B1_o , \t/a/aluin/sel0_b13/B0 , \t/a/aluin/sel0_b13/B1 );
  or \t/a/aluin/sel0_b13/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b13/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b13/B2 , \t/a/aluin/sel0_b13/B3 );
  or \t/a/aluin/sel0_b13/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [13], \t/a/aluin/sel0_b13/or_B0_B1_o , \t/a/aluin/sel0_b13/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b14/and_b0_0  (\t/a/aluin/sel0_b14/B0 , \t/a/aluin/o_A1 [14], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b14/and_b0_1  (\t/a/aluin/sel0_b14/B1 , \t/a/EX_memstraddr [14], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b14/and_b0_2  (\t/a/aluin/sel0_b14/B2 , \t/a/EX_memstraddr [14], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b14/and_b0_3  (\t/a/aluin/sel0_b14/B3 , \t/a/EX_memstraddr [14], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b14/or_B0_B1  (\t/a/aluin/sel0_b14/or_B0_B1_o , \t/a/aluin/sel0_b14/B0 , \t/a/aluin/sel0_b14/B1 );
  or \t/a/aluin/sel0_b14/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b14/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b14/B2 , \t/a/aluin/sel0_b14/B3 );
  or \t/a/aluin/sel0_b14/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [14], \t/a/aluin/sel0_b14/or_B0_B1_o , \t/a/aluin/sel0_b14/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b15/and_b0_0  (\t/a/aluin/sel0_b15/B0 , \t/a/aluin/o_A1 [15], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b15/and_b0_1  (\t/a/aluin/sel0_b15/B1 , \t/a/EX_memstraddr [15], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b15/and_b0_2  (\t/a/aluin/sel0_b15/B2 , \t/a/EX_memstraddr [15], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b15/and_b0_3  (\t/a/aluin/sel0_b15/B3 , \t/a/EX_memstraddr [15], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b15/or_B0_B1  (\t/a/aluin/sel0_b15/or_B0_B1_o , \t/a/aluin/sel0_b15/B0 , \t/a/aluin/sel0_b15/B1 );
  or \t/a/aluin/sel0_b15/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b15/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b15/B2 , \t/a/aluin/sel0_b15/B3 );
  or \t/a/aluin/sel0_b15/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [15], \t/a/aluin/sel0_b15/or_B0_B1_o , \t/a/aluin/sel0_b15/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b16/and_b0_0  (\t/a/aluin/sel0_b16/B0 , \t/a/aluin/o_A1 [16], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b16/and_b0_1  (\t/a/aluin/sel0_b16/B1 , \t/a/EX_memstraddr [16], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b16/and_b0_2  (\t/a/aluin/sel0_b16/B2 , \t/a/EX_memstraddr [16], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b16/and_b0_3  (\t/a/aluin/sel0_b16/B3 , \t/a/EX_memstraddr [16], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b16/or_B0_B1  (\t/a/aluin/sel0_b16/or_B0_B1_o , \t/a/aluin/sel0_b16/B0 , \t/a/aluin/sel0_b16/B1 );
  or \t/a/aluin/sel0_b16/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b16/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b16/B2 , \t/a/aluin/sel0_b16/B3 );
  or \t/a/aluin/sel0_b16/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [16], \t/a/aluin/sel0_b16/or_B0_B1_o , \t/a/aluin/sel0_b16/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b17/and_b0_0  (\t/a/aluin/sel0_b17/B0 , \t/a/aluin/o_A1 [17], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b17/and_b0_1  (\t/a/aluin/sel0_b17/B1 , \t/a/EX_memstraddr [17], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b17/and_b0_2  (\t/a/aluin/sel0_b17/B2 , \t/a/EX_memstraddr [17], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b17/and_b0_3  (\t/a/aluin/sel0_b17/B3 , \t/a/EX_memstraddr [17], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b17/or_B0_B1  (\t/a/aluin/sel0_b17/or_B0_B1_o , \t/a/aluin/sel0_b17/B0 , \t/a/aluin/sel0_b17/B1 );
  or \t/a/aluin/sel0_b17/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b17/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b17/B2 , \t/a/aluin/sel0_b17/B3 );
  or \t/a/aluin/sel0_b17/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [17], \t/a/aluin/sel0_b17/or_B0_B1_o , \t/a/aluin/sel0_b17/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b18/and_b0_0  (\t/a/aluin/sel0_b18/B0 , \t/a/aluin/o_A1 [18], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b18/and_b0_1  (\t/a/aluin/sel0_b18/B1 , \t/a/EX_memstraddr [18], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b18/and_b0_2  (\t/a/aluin/sel0_b18/B2 , \t/a/EX_memstraddr [18], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b18/and_b0_3  (\t/a/aluin/sel0_b18/B3 , \t/a/EX_memstraddr [18], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b18/or_B0_B1  (\t/a/aluin/sel0_b18/or_B0_B1_o , \t/a/aluin/sel0_b18/B0 , \t/a/aluin/sel0_b18/B1 );
  or \t/a/aluin/sel0_b18/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b18/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b18/B2 , \t/a/aluin/sel0_b18/B3 );
  or \t/a/aluin/sel0_b18/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [18], \t/a/aluin/sel0_b18/or_B0_B1_o , \t/a/aluin/sel0_b18/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b19/and_b0_0  (\t/a/aluin/sel0_b19/B0 , \t/a/aluin/o_A1 [19], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b19/and_b0_1  (\t/a/aluin/sel0_b19/B1 , \t/a/EX_memstraddr [19], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b19/and_b0_2  (\t/a/aluin/sel0_b19/B2 , \t/a/EX_memstraddr [19], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b19/and_b0_3  (\t/a/aluin/sel0_b19/B3 , \t/a/EX_memstraddr [19], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b19/or_B0_B1  (\t/a/aluin/sel0_b19/or_B0_B1_o , \t/a/aluin/sel0_b19/B0 , \t/a/aluin/sel0_b19/B1 );
  or \t/a/aluin/sel0_b19/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b19/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b19/B2 , \t/a/aluin/sel0_b19/B3 );
  or \t/a/aluin/sel0_b19/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [19], \t/a/aluin/sel0_b19/or_B0_B1_o , \t/a/aluin/sel0_b19/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b2/and_b0_0  (\t/a/aluin/sel0_b2/B0 , \t/a/aluin/o_A1 [2], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b2/and_b0_1  (\t/a/aluin/sel0_b2/B1 , \t/a/EX_memstraddr [2], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b2/and_b0_2  (\t/a/aluin/sel0_b2/B2 , \t/a/EX_memstraddr [2], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b2/and_b0_3  (\t/a/aluin/sel0_b2/B3 , \t/a/EX_memstraddr [2], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b2/or_B0_B1  (\t/a/aluin/sel0_b2/or_B0_B1_o , \t/a/aluin/sel0_b2/B0 , \t/a/aluin/sel0_b2/B1 );
  or \t/a/aluin/sel0_b2/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b2/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b2/B2 , \t/a/aluin/sel0_b2/B3 );
  or \t/a/aluin/sel0_b2/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [2], \t/a/aluin/sel0_b2/or_B0_B1_o , \t/a/aluin/sel0_b2/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b20/and_b0_0  (\t/a/aluin/sel0_b20/B0 , \t/a/aluin/o_A1 [20], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b20/and_b0_1  (\t/a/aluin/sel0_b20/B1 , \t/a/EX_memstraddr [20], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b20/and_b0_2  (\t/a/aluin/sel0_b20/B2 , \t/a/EX_memstraddr [20], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b20/and_b0_3  (\t/a/aluin/sel0_b20/B3 , \t/a/EX_memstraddr [20], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b20/or_B0_B1  (\t/a/aluin/sel0_b20/or_B0_B1_o , \t/a/aluin/sel0_b20/B0 , \t/a/aluin/sel0_b20/B1 );
  or \t/a/aluin/sel0_b20/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b20/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b20/B2 , \t/a/aluin/sel0_b20/B3 );
  or \t/a/aluin/sel0_b20/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [20], \t/a/aluin/sel0_b20/or_B0_B1_o , \t/a/aluin/sel0_b20/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b21/and_b0_0  (\t/a/aluin/sel0_b21/B0 , \t/a/aluin/o_A1 [21], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b21/and_b0_1  (\t/a/aluin/sel0_b21/B1 , \t/a/EX_memstraddr [21], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b21/and_b0_2  (\t/a/aluin/sel0_b21/B2 , \t/a/EX_memstraddr [21], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b21/and_b0_3  (\t/a/aluin/sel0_b21/B3 , \t/a/EX_memstraddr [21], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b21/or_B0_B1  (\t/a/aluin/sel0_b21/or_B0_B1_o , \t/a/aluin/sel0_b21/B0 , \t/a/aluin/sel0_b21/B1 );
  or \t/a/aluin/sel0_b21/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b21/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b21/B2 , \t/a/aluin/sel0_b21/B3 );
  or \t/a/aluin/sel0_b21/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [21], \t/a/aluin/sel0_b21/or_B0_B1_o , \t/a/aluin/sel0_b21/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b22/and_b0_0  (\t/a/aluin/sel0_b22/B0 , \t/a/aluin/o_A1 [22], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b22/and_b0_1  (\t/a/aluin/sel0_b22/B1 , \t/a/EX_memstraddr [22], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b22/and_b0_2  (\t/a/aluin/sel0_b22/B2 , \t/a/EX_memstraddr [22], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b22/and_b0_3  (\t/a/aluin/sel0_b22/B3 , \t/a/EX_memstraddr [22], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b22/or_B0_B1  (\t/a/aluin/sel0_b22/or_B0_B1_o , \t/a/aluin/sel0_b22/B0 , \t/a/aluin/sel0_b22/B1 );
  or \t/a/aluin/sel0_b22/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b22/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b22/B2 , \t/a/aluin/sel0_b22/B3 );
  or \t/a/aluin/sel0_b22/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [22], \t/a/aluin/sel0_b22/or_B0_B1_o , \t/a/aluin/sel0_b22/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b23/and_b0_0  (\t/a/aluin/sel0_b23/B0 , \t/a/aluin/o_A1 [23], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b23/and_b0_1  (\t/a/aluin/sel0_b23/B1 , \t/a/EX_memstraddr [23], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b23/and_b0_2  (\t/a/aluin/sel0_b23/B2 , \t/a/EX_memstraddr [23], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b23/and_b0_3  (\t/a/aluin/sel0_b23/B3 , \t/a/EX_memstraddr [23], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b23/or_B0_B1  (\t/a/aluin/sel0_b23/or_B0_B1_o , \t/a/aluin/sel0_b23/B0 , \t/a/aluin/sel0_b23/B1 );
  or \t/a/aluin/sel0_b23/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b23/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b23/B2 , \t/a/aluin/sel0_b23/B3 );
  or \t/a/aluin/sel0_b23/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [23], \t/a/aluin/sel0_b23/or_B0_B1_o , \t/a/aluin/sel0_b23/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b24/and_b0_0  (\t/a/aluin/sel0_b24/B0 , \t/a/aluin/o_A1 [24], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b24/and_b0_1  (\t/a/aluin/sel0_b24/B1 , \t/a/EX_memstraddr [24], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b24/and_b0_2  (\t/a/aluin/sel0_b24/B2 , \t/a/EX_memstraddr [24], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b24/and_b0_3  (\t/a/aluin/sel0_b24/B3 , \t/a/EX_memstraddr [24], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b24/or_B0_B1  (\t/a/aluin/sel0_b24/or_B0_B1_o , \t/a/aluin/sel0_b24/B0 , \t/a/aluin/sel0_b24/B1 );
  or \t/a/aluin/sel0_b24/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b24/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b24/B2 , \t/a/aluin/sel0_b24/B3 );
  or \t/a/aluin/sel0_b24/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [24], \t/a/aluin/sel0_b24/or_B0_B1_o , \t/a/aluin/sel0_b24/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b25/and_b0_0  (\t/a/aluin/sel0_b25/B0 , \t/a/aluin/o_A1 [25], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b25/and_b0_1  (\t/a/aluin/sel0_b25/B1 , \t/a/EX_memstraddr [25], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b25/and_b0_2  (\t/a/aluin/sel0_b25/B2 , \t/a/EX_memstraddr [25], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b25/and_b0_3  (\t/a/aluin/sel0_b25/B3 , \t/a/EX_memstraddr [25], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b25/or_B0_B1  (\t/a/aluin/sel0_b25/or_B0_B1_o , \t/a/aluin/sel0_b25/B0 , \t/a/aluin/sel0_b25/B1 );
  or \t/a/aluin/sel0_b25/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b25/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b25/B2 , \t/a/aluin/sel0_b25/B3 );
  or \t/a/aluin/sel0_b25/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [25], \t/a/aluin/sel0_b25/or_B0_B1_o , \t/a/aluin/sel0_b25/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b26/and_b0_0  (\t/a/aluin/sel0_b26/B0 , \t/a/aluin/o_A1 [26], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b26/and_b0_1  (\t/a/aluin/sel0_b26/B1 , \t/a/EX_memstraddr [26], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b26/and_b0_2  (\t/a/aluin/sel0_b26/B2 , \t/a/EX_memstraddr [26], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b26/and_b0_3  (\t/a/aluin/sel0_b26/B3 , \t/a/EX_memstraddr [26], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b26/or_B0_B1  (\t/a/aluin/sel0_b26/or_B0_B1_o , \t/a/aluin/sel0_b26/B0 , \t/a/aluin/sel0_b26/B1 );
  or \t/a/aluin/sel0_b26/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b26/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b26/B2 , \t/a/aluin/sel0_b26/B3 );
  or \t/a/aluin/sel0_b26/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [26], \t/a/aluin/sel0_b26/or_B0_B1_o , \t/a/aluin/sel0_b26/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b27/and_b0_0  (\t/a/aluin/sel0_b27/B0 , \t/a/aluin/o_A1 [27], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b27/and_b0_1  (\t/a/aluin/sel0_b27/B1 , \t/a/EX_memstraddr [27], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b27/and_b0_2  (\t/a/aluin/sel0_b27/B2 , \t/a/EX_memstraddr [27], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b27/and_b0_3  (\t/a/aluin/sel0_b27/B3 , \t/a/EX_memstraddr [27], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b27/or_B0_B1  (\t/a/aluin/sel0_b27/or_B0_B1_o , \t/a/aluin/sel0_b27/B0 , \t/a/aluin/sel0_b27/B1 );
  or \t/a/aluin/sel0_b27/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b27/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b27/B2 , \t/a/aluin/sel0_b27/B3 );
  or \t/a/aluin/sel0_b27/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [27], \t/a/aluin/sel0_b27/or_B0_B1_o , \t/a/aluin/sel0_b27/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b28/and_b0_0  (\t/a/aluin/sel0_b28/B0 , \t/a/aluin/o_A1 [28], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b28/and_b0_1  (\t/a/aluin/sel0_b28/B1 , \t/a/EX_memstraddr [28], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b28/and_b0_2  (\t/a/aluin/sel0_b28/B2 , \t/a/EX_memstraddr [28], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b28/and_b0_3  (\t/a/aluin/sel0_b28/B3 , \t/a/EX_memstraddr [28], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b28/or_B0_B1  (\t/a/aluin/sel0_b28/or_B0_B1_o , \t/a/aluin/sel0_b28/B0 , \t/a/aluin/sel0_b28/B1 );
  or \t/a/aluin/sel0_b28/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b28/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b28/B2 , \t/a/aluin/sel0_b28/B3 );
  or \t/a/aluin/sel0_b28/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [28], \t/a/aluin/sel0_b28/or_B0_B1_o , \t/a/aluin/sel0_b28/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b29/and_b0_0  (\t/a/aluin/sel0_b29/B0 , \t/a/aluin/o_A1 [29], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b29/and_b0_1  (\t/a/aluin/sel0_b29/B1 , \t/a/EX_memstraddr [29], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b29/and_b0_2  (\t/a/aluin/sel0_b29/B2 , \t/a/EX_memstraddr [29], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b29/and_b0_3  (\t/a/aluin/sel0_b29/B3 , \t/a/EX_memstraddr [29], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b29/or_B0_B1  (\t/a/aluin/sel0_b29/or_B0_B1_o , \t/a/aluin/sel0_b29/B0 , \t/a/aluin/sel0_b29/B1 );
  or \t/a/aluin/sel0_b29/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b29/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b29/B2 , \t/a/aluin/sel0_b29/B3 );
  or \t/a/aluin/sel0_b29/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [29], \t/a/aluin/sel0_b29/or_B0_B1_o , \t/a/aluin/sel0_b29/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b3/and_b0_0  (\t/a/aluin/sel0_b3/B0 , \t/a/aluin/o_A1 [3], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b3/and_b0_1  (\t/a/aluin/sel0_b3/B1 , \t/a/EX_memstraddr [3], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b3/and_b0_2  (\t/a/aluin/sel0_b3/B2 , \t/a/EX_memstraddr [3], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b3/and_b0_3  (\t/a/aluin/sel0_b3/B3 , \t/a/EX_memstraddr [3], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b3/or_B0_B1  (\t/a/aluin/sel0_b3/or_B0_B1_o , \t/a/aluin/sel0_b3/B0 , \t/a/aluin/sel0_b3/B1 );
  or \t/a/aluin/sel0_b3/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b3/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b3/B2 , \t/a/aluin/sel0_b3/B3 );
  or \t/a/aluin/sel0_b3/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [3], \t/a/aluin/sel0_b3/or_B0_B1_o , \t/a/aluin/sel0_b3/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b30/and_b0_0  (\t/a/aluin/sel0_b30/B0 , \t/a/aluin/o_A1 [30], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b30/and_b0_1  (\t/a/aluin/sel0_b30/B1 , \t/a/EX_memstraddr [30], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b30/and_b0_2  (\t/a/aluin/sel0_b30/B2 , \t/a/EX_memstraddr [30], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b30/and_b0_3  (\t/a/aluin/sel0_b30/B3 , \t/a/EX_memstraddr [30], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b30/or_B0_B1  (\t/a/aluin/sel0_b30/or_B0_B1_o , \t/a/aluin/sel0_b30/B0 , \t/a/aluin/sel0_b30/B1 );
  or \t/a/aluin/sel0_b30/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b30/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b30/B2 , \t/a/aluin/sel0_b30/B3 );
  or \t/a/aluin/sel0_b30/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [30], \t/a/aluin/sel0_b30/or_B0_B1_o , \t/a/aluin/sel0_b30/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b31/and_b0_0  (\t/a/aluin/sel0_b31/B0 , \t/a/aluin/o_A1 [31], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b31/and_b0_1  (\t/a/aluin/sel0_b31/B1 , \t/a/EX_memstraddr [31], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b31/and_b0_2  (\t/a/aluin/sel0_b31/B2 , \t/a/EX_memstraddr [31], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b31/and_b0_3  (\t/a/aluin/sel0_b31/B3 , \t/a/EX_memstraddr [31], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b31/or_B0_B1  (\t/a/aluin/sel0_b31/or_B0_B1_o , \t/a/aluin/sel0_b31/B0 , \t/a/aluin/sel0_b31/B1 );
  or \t/a/aluin/sel0_b31/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b31/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b31/B2 , \t/a/aluin/sel0_b31/B3 );
  or \t/a/aluin/sel0_b31/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [31], \t/a/aluin/sel0_b31/or_B0_B1_o , \t/a/aluin/sel0_b31/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b4/and_b0_0  (\t/a/aluin/sel0_b4/B0 , \t/a/aluin/o_A1 [4], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b4/and_b0_1  (\t/a/aluin/sel0_b4/B1 , \t/a/EX_memstraddr [4], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b4/and_b0_2  (\t/a/aluin/sel0_b4/B2 , \t/a/EX_memstraddr [4], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b4/and_b0_3  (\t/a/aluin/sel0_b4/B3 , \t/a/EX_memstraddr [4], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b4/or_B0_B1  (\t/a/aluin/sel0_b4/or_B0_B1_o , \t/a/aluin/sel0_b4/B0 , \t/a/aluin/sel0_b4/B1 );
  or \t/a/aluin/sel0_b4/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b4/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b4/B2 , \t/a/aluin/sel0_b4/B3 );
  or \t/a/aluin/sel0_b4/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [4], \t/a/aluin/sel0_b4/or_B0_B1_o , \t/a/aluin/sel0_b4/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b5/and_b0_0  (\t/a/aluin/sel0_b5/B0 , \t/a/aluin/o_A1 [5], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b5/and_b0_1  (\t/a/aluin/sel0_b5/B1 , \t/a/EX_memstraddr [5], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b5/and_b0_2  (\t/a/aluin/sel0_b5/B2 , \t/a/EX_memstraddr [5], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b5/and_b0_3  (\t/a/aluin/sel0_b5/B3 , \t/a/EX_memstraddr [5], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b5/or_B0_B1  (\t/a/aluin/sel0_b5/or_B0_B1_o , \t/a/aluin/sel0_b5/B0 , \t/a/aluin/sel0_b5/B1 );
  or \t/a/aluin/sel0_b5/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b5/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b5/B2 , \t/a/aluin/sel0_b5/B3 );
  or \t/a/aluin/sel0_b5/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [5], \t/a/aluin/sel0_b5/or_B0_B1_o , \t/a/aluin/sel0_b5/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b6/and_b0_0  (\t/a/aluin/sel0_b6/B0 , \t/a/aluin/o_A1 [6], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b6/and_b0_1  (\t/a/aluin/sel0_b6/B1 , \t/a/EX_memstraddr [6], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b6/and_b0_2  (\t/a/aluin/sel0_b6/B2 , \t/a/EX_memstraddr [6], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b6/and_b0_3  (\t/a/aluin/sel0_b6/B3 , \t/a/EX_memstraddr [6], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b6/or_B0_B1  (\t/a/aluin/sel0_b6/or_B0_B1_o , \t/a/aluin/sel0_b6/B0 , \t/a/aluin/sel0_b6/B1 );
  or \t/a/aluin/sel0_b6/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b6/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b6/B2 , \t/a/aluin/sel0_b6/B3 );
  or \t/a/aluin/sel0_b6/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [6], \t/a/aluin/sel0_b6/or_B0_B1_o , \t/a/aluin/sel0_b6/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b7/and_b0_0  (\t/a/aluin/sel0_b7/B0 , \t/a/aluin/o_A1 [7], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b7/and_b0_1  (\t/a/aluin/sel0_b7/B1 , \t/a/EX_memstraddr [7], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b7/and_b0_2  (\t/a/aluin/sel0_b7/B2 , \t/a/EX_memstraddr [7], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b7/and_b0_3  (\t/a/aluin/sel0_b7/B3 , \t/a/EX_memstraddr [7], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b7/or_B0_B1  (\t/a/aluin/sel0_b7/or_B0_B1_o , \t/a/aluin/sel0_b7/B0 , \t/a/aluin/sel0_b7/B1 );
  or \t/a/aluin/sel0_b7/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b7/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b7/B2 , \t/a/aluin/sel0_b7/B3 );
  or \t/a/aluin/sel0_b7/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [7], \t/a/aluin/sel0_b7/or_B0_B1_o , \t/a/aluin/sel0_b7/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b8/and_b0_0  (\t/a/aluin/sel0_b8/B0 , \t/a/aluin/o_A1 [8], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b8/and_b0_1  (\t/a/aluin/sel0_b8/B1 , \t/a/EX_memstraddr [8], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b8/and_b0_2  (\t/a/aluin/sel0_b8/B2 , \t/a/EX_memstraddr [8], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b8/and_b0_3  (\t/a/aluin/sel0_b8/B3 , \t/a/EX_memstraddr [8], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b8/or_B0_B1  (\t/a/aluin/sel0_b8/or_B0_B1_o , \t/a/aluin/sel0_b8/B0 , \t/a/aluin/sel0_b8/B1 );
  or \t/a/aluin/sel0_b8/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b8/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b8/B2 , \t/a/aluin/sel0_b8/B3 );
  or \t/a/aluin/sel0_b8/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [8], \t/a/aluin/sel0_b8/or_B0_B1_o , \t/a/aluin/sel0_b8/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel0_b9/and_b0_0  (\t/a/aluin/sel0_b9/B0 , \t/a/aluin/o_A1 [9], \t/a/aluin/n5 );
  and \t/a/aluin/sel0_b9/and_b0_1  (\t/a/aluin/sel0_b9/B1 , \t/a/EX_memstraddr [9], \t/a/aluin/n4 );
  and \t/a/aluin/sel0_b9/and_b0_2  (\t/a/aluin/sel0_b9/B2 , \t/a/EX_memstraddr [9], \t/a/aluin/n3 );
  and \t/a/aluin/sel0_b9/and_b0_3  (\t/a/aluin/sel0_b9/B3 , \t/a/EX_memstraddr [9], \t/a/aluin/n2 );
  or \t/a/aluin/sel0_b9/or_B0_B1  (\t/a/aluin/sel0_b9/or_B0_B1_o , \t/a/aluin/sel0_b9/B0 , \t/a/aluin/sel0_b9/B1 );
  or \t/a/aluin/sel0_b9/or_B2_or_B3_B4_o  (\t/a/aluin/sel0_b9/or_B2_or_B3_B4_o_o , \t/a/aluin/sel0_b9/B2 , \t/a/aluin/sel0_b9/B3 );
  or \t/a/aluin/sel0_b9/or_or_B0_B1_o_or_B2_  (\t/a/EX_A [9], \t/a/aluin/sel0_b9/or_B0_B1_o , \t/a/aluin/sel0_b9/or_B2_or_B3_B4_o_o );
  and \t/a/aluin/sel1_b0/and_b0_6  (\t/a/aluin/sel1_b0/B6 , \t/a/EX_rs2 [0], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b0/and_b0_7  (\t/a/aluin/sel1_b0/B7 , \t/a/EX_rd [0], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b0/and_b0_8  (\t/a/aluin/sel1_b0/B8 , \t/a/EX_rs2 [0], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b0/and_b0_9  (\t/a/aluin/sel1_b0/B9 , \t/a/aluin/o_B1 [0], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b0/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b0/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b0/B7 , \t/a/aluin/sel1_b0/or_B8_B9_o );
  or \t/a/aluin/sel1_b0/or_B8_B9  (\t/a/aluin/sel1_b0/or_B8_B9_o , \t/a/aluin/sel1_b0/B8 , \t/a/aluin/sel1_b0/B9 );
  or \t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b0/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b0/B6 , \t/a/aluin/sel1_b0/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b1/and_b0_6  (\t/a/aluin/sel1_b1/B6 , \t/a/EX_rs2 [1], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b1/and_b0_7  (\t/a/aluin/sel1_b1/B7 , \t/a/EX_rd [1], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b1/and_b0_8  (\t/a/aluin/sel1_b1/B8 , \t/a/EX_rs2 [1], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b1/and_b0_9  (\t/a/aluin/sel1_b1/B9 , \t/a/aluin/o_B1 [1], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b1/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b1/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b1/B7 , \t/a/aluin/sel1_b1/or_B8_B9_o );
  or \t/a/aluin/sel1_b1/or_B8_B9  (\t/a/aluin/sel1_b1/or_B8_B9_o , \t/a/aluin/sel1_b1/B8 , \t/a/aluin/sel1_b1/B9 );
  or \t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b1/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b1/B6 , \t/a/aluin/sel1_b1/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b10/and_b0_6  (\t/a/aluin/sel1_b10/B6 , \t/a/aluin/n9 [5], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b10/and_b0_7  (\t/a/aluin/sel1_b10/B7 , \t/a/EX_fun7 [5], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b10/and_b0_8  (\t/a/aluin/sel1_b10/B8 , \t/a/EX_fun7 [5], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b10/and_b0_9  (\t/a/aluin/sel1_b10/B9 , \t/a/aluin/o_B1 [10], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b10/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b10/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b10/B7 , \t/a/aluin/sel1_b10/or_B8_B9_o );
  or \t/a/aluin/sel1_b10/or_B8_B9  (\t/a/aluin/sel1_b10/or_B8_B9_o , \t/a/aluin/sel1_b10/B8 , \t/a/aluin/sel1_b10/B9 );
  or \t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b10/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b10/B6 , \t/a/aluin/sel1_b10/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b11/and_b0_6  (\t/a/aluin/sel1_b11/B6 , \t/a/aluin/n9 [6], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b11/and_b0_7  (\t/a/aluin/sel1_b11/B7 , \t/a/EX_fun7 [6], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b11/and_b0_8  (\t/a/aluin/sel1_b11/B8 , \t/a/EX_fun7 [6], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b11/and_b0_9  (\t/a/aluin/sel1_b11/B9 , \t/a/aluin/o_B1 [11], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b11/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b11/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b11/or_B8_B9_o );
  or \t/a/aluin/sel1_b11/or_B8_B9  (\t/a/aluin/sel1_b11/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b11/B9 );
  or \t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b11/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b11/B6 , \t/a/aluin/sel1_b11/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b12/and_b0_2  (\t/a/aluin/sel1_b12/B2 , \t/a/EX_fun3 [0], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b12/and_b0_3  (\t/a/aluin/sel1_b12/B3 , \t/a/EX_fun3 [0], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b12/and_b0_9  (\t/a/aluin/sel1_b12/B9 , \t/a/aluin/o_B1 [12], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b12/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b12/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b12/B2 , \t/a/aluin/sel1_b12/B3 );
  or \t/a/aluin/sel1_b12/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b12/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b12/or_B8_B9_o );
  or \t/a/aluin/sel1_b12/or_B8_B9  (\t/a/aluin/sel1_b12/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b12/B9 );
  or \t/a/aluin/sel1_b12/or_or_or_B0_B1_o_or_  (\t/a/EX_B [12], \t/a/aluin/sel1_b12/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b12/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b13/and_b0_2  (\t/a/aluin/sel1_b13/B2 , \t/a/EX_fun3 [1], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b13/and_b0_3  (\t/a/aluin/sel1_b13/B3 , \t/a/EX_fun3 [1], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b13/and_b0_9  (\t/a/aluin/sel1_b13/B9 , \t/a/aluin/o_B1 [13], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b13/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b13/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b13/B2 , \t/a/aluin/sel1_b13/B3 );
  or \t/a/aluin/sel1_b13/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b13/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b13/or_B8_B9_o );
  or \t/a/aluin/sel1_b13/or_B8_B9  (\t/a/aluin/sel1_b13/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b13/B9 );
  or \t/a/aluin/sel1_b13/or_or_or_B0_B1_o_or_  (\t/a/EX_B [13], \t/a/aluin/sel1_b13/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b13/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b14/and_b0_2  (\t/a/aluin/sel1_b14/B2 , \t/a/EX_fun3 [2], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b14/and_b0_3  (\t/a/aluin/sel1_b14/B3 , \t/a/EX_fun3 [2], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b14/and_b0_9  (\t/a/aluin/sel1_b14/B9 , \t/a/aluin/o_B1 [14], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b14/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b14/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b14/B2 , \t/a/aluin/sel1_b14/B3 );
  or \t/a/aluin/sel1_b14/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b14/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b14/or_B8_B9_o );
  or \t/a/aluin/sel1_b14/or_B8_B9  (\t/a/aluin/sel1_b14/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b14/B9 );
  or \t/a/aluin/sel1_b14/or_or_or_B0_B1_o_or_  (\t/a/EX_B [14], \t/a/aluin/sel1_b14/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b14/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b15/and_b0_2  (\t/a/aluin/sel1_b15/B2 , \t/a/EX_rs1 [0], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b15/and_b0_3  (\t/a/aluin/sel1_b15/B3 , \t/a/EX_rs1 [0], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b15/and_b0_9  (\t/a/aluin/sel1_b15/B9 , \t/a/aluin/o_B1 [15], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b15/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b15/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b15/B2 , \t/a/aluin/sel1_b15/B3 );
  or \t/a/aluin/sel1_b15/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b15/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b15/or_B8_B9_o );
  or \t/a/aluin/sel1_b15/or_B8_B9  (\t/a/aluin/sel1_b15/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b15/B9 );
  or \t/a/aluin/sel1_b15/or_or_or_B0_B1_o_or_  (\t/a/EX_B [15], \t/a/aluin/sel1_b15/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b15/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b16/and_b0_2  (\t/a/aluin/sel1_b16/B2 , \t/a/EX_rs1 [1], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b16/and_b0_3  (\t/a/aluin/sel1_b16/B3 , \t/a/EX_rs1 [1], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b16/and_b0_9  (\t/a/aluin/sel1_b16/B9 , \t/a/aluin/o_B1 [16], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b16/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b16/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b16/B2 , \t/a/aluin/sel1_b16/B3 );
  or \t/a/aluin/sel1_b16/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b16/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b16/or_B8_B9_o );
  or \t/a/aluin/sel1_b16/or_B8_B9  (\t/a/aluin/sel1_b16/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b16/B9 );
  or \t/a/aluin/sel1_b16/or_or_or_B0_B1_o_or_  (\t/a/EX_B [16], \t/a/aluin/sel1_b16/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b16/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b17/and_b0_2  (\t/a/aluin/sel1_b17/B2 , \t/a/EX_rs1 [2], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b17/and_b0_3  (\t/a/aluin/sel1_b17/B3 , \t/a/EX_rs1 [2], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b17/and_b0_9  (\t/a/aluin/sel1_b17/B9 , \t/a/aluin/o_B1 [17], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b17/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b17/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b17/B2 , \t/a/aluin/sel1_b17/B3 );
  or \t/a/aluin/sel1_b17/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b17/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b17/or_B8_B9_o );
  or \t/a/aluin/sel1_b17/or_B8_B9  (\t/a/aluin/sel1_b17/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b17/B9 );
  or \t/a/aluin/sel1_b17/or_or_or_B0_B1_o_or_  (\t/a/EX_B [17], \t/a/aluin/sel1_b17/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b17/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b18/and_b0_2  (\t/a/aluin/sel1_b18/B2 , \t/a/EX_rs1 [3], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b18/and_b0_3  (\t/a/aluin/sel1_b18/B3 , \t/a/EX_rs1 [3], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b18/and_b0_9  (\t/a/aluin/sel1_b18/B9 , \t/a/aluin/o_B1 [18], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b18/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b18/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b18/B2 , \t/a/aluin/sel1_b18/B3 );
  or \t/a/aluin/sel1_b18/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b18/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b18/or_B8_B9_o );
  or \t/a/aluin/sel1_b18/or_B8_B9  (\t/a/aluin/sel1_b18/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b18/B9 );
  or \t/a/aluin/sel1_b18/or_or_or_B0_B1_o_or_  (\t/a/EX_B [18], \t/a/aluin/sel1_b18/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b18/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b19/and_b0_2  (\t/a/aluin/sel1_b19/B2 , \t/a/EX_rs1 [4], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b19/and_b0_3  (\t/a/aluin/sel1_b19/B3 , \t/a/EX_rs1 [4], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b19/and_b0_9  (\t/a/aluin/sel1_b19/B9 , \t/a/aluin/o_B1 [19], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b19/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b19/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b19/B2 , \t/a/aluin/sel1_b19/B3 );
  or \t/a/aluin/sel1_b19/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b19/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b19/or_B8_B9_o );
  or \t/a/aluin/sel1_b19/or_B8_B9  (\t/a/aluin/sel1_b19/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b19/B9 );
  or \t/a/aluin/sel1_b19/or_or_or_B0_B1_o_or_  (\t/a/EX_B [19], \t/a/aluin/sel1_b19/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b19/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b2/and_b0_6  (\t/a/aluin/sel1_b2/B6 , \t/a/EX_rs2 [2], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b2/and_b0_7  (\t/a/aluin/sel1_b2/B7 , \t/a/EX_rd [2], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b2/and_b0_8  (\t/a/aluin/sel1_b2/B8 , \t/a/EX_rs2 [2], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b2/and_b0_9  (\t/a/aluin/sel1_b2/B9 , \t/a/aluin/o_B1 [2], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b2/or_B5_B6  (\t/a/aluin/sel1_b2/or_B5_B6_o , \t/a/aluin/n2 , \t/a/aluin/sel1_b2/B6 );
  or \t/a/aluin/sel1_b2/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b2/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b2/B7 , \t/a/aluin/sel1_b2/or_B8_B9_o );
  or \t/a/aluin/sel1_b2/or_B8_B9  (\t/a/aluin/sel1_b2/or_B8_B9_o , \t/a/aluin/sel1_b2/B8 , \t/a/aluin/sel1_b2/B9 );
  or \t/a/aluin/sel1_b2/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b2/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b2/or_B5_B6_o , \t/a/aluin/sel1_b2/or_B7_or_B8_B9_o_o );
  or \t/a/aluin/sel1_b2/or_or_or_B0_B1_o_or_  (\t/a/EX_B [2], \t/a/aluin/n3 , \t/a/aluin/sel1_b2/or_or_B5_B6_o_or_B7__o );
  and \t/a/aluin/sel1_b20/and_b0_2  (\t/a/aluin/sel1_b20/B2 , \t/a/EX_rs2 [0], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b20/and_b0_3  (\t/a/aluin/sel1_b20/B3 , \t/a/EX_rs2 [0], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b20/and_b0_9  (\t/a/aluin/sel1_b20/B9 , \t/a/aluin/o_B1 [20], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b20/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b20/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b20/B2 , \t/a/aluin/sel1_b20/B3 );
  or \t/a/aluin/sel1_b20/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b20/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b20/or_B8_B9_o );
  or \t/a/aluin/sel1_b20/or_B8_B9  (\t/a/aluin/sel1_b20/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b20/B9 );
  or \t/a/aluin/sel1_b20/or_or_or_B0_B1_o_or_  (\t/a/EX_B [20], \t/a/aluin/sel1_b20/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b20/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b21/and_b0_2  (\t/a/aluin/sel1_b21/B2 , \t/a/EX_rs2 [1], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b21/and_b0_3  (\t/a/aluin/sel1_b21/B3 , \t/a/EX_rs2 [1], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b21/and_b0_9  (\t/a/aluin/sel1_b21/B9 , \t/a/aluin/o_B1 [21], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b21/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b21/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b21/B2 , \t/a/aluin/sel1_b21/B3 );
  or \t/a/aluin/sel1_b21/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b21/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b21/or_B8_B9_o );
  or \t/a/aluin/sel1_b21/or_B8_B9  (\t/a/aluin/sel1_b21/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b21/B9 );
  or \t/a/aluin/sel1_b21/or_or_or_B0_B1_o_or_  (\t/a/EX_B [21], \t/a/aluin/sel1_b21/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b21/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b22/and_b0_2  (\t/a/aluin/sel1_b22/B2 , \t/a/EX_rs2 [2], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b22/and_b0_3  (\t/a/aluin/sel1_b22/B3 , \t/a/EX_rs2 [2], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b22/and_b0_9  (\t/a/aluin/sel1_b22/B9 , \t/a/aluin/o_B1 [22], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b22/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b22/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b22/B2 , \t/a/aluin/sel1_b22/B3 );
  or \t/a/aluin/sel1_b22/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b22/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b22/or_B8_B9_o );
  or \t/a/aluin/sel1_b22/or_B8_B9  (\t/a/aluin/sel1_b22/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b22/B9 );
  or \t/a/aluin/sel1_b22/or_or_or_B0_B1_o_or_  (\t/a/EX_B [22], \t/a/aluin/sel1_b22/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b22/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b23/and_b0_2  (\t/a/aluin/sel1_b23/B2 , \t/a/EX_rs2 [3], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b23/and_b0_3  (\t/a/aluin/sel1_b23/B3 , \t/a/EX_rs2 [3], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b23/and_b0_9  (\t/a/aluin/sel1_b23/B9 , \t/a/aluin/o_B1 [23], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b23/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b23/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b23/B2 , \t/a/aluin/sel1_b23/B3 );
  or \t/a/aluin/sel1_b23/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b23/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b23/or_B8_B9_o );
  or \t/a/aluin/sel1_b23/or_B8_B9  (\t/a/aluin/sel1_b23/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b23/B9 );
  or \t/a/aluin/sel1_b23/or_or_or_B0_B1_o_or_  (\t/a/EX_B [23], \t/a/aluin/sel1_b23/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b23/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b24/and_b0_2  (\t/a/aluin/sel1_b24/B2 , \t/a/EX_rs2 [4], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b24/and_b0_3  (\t/a/aluin/sel1_b24/B3 , \t/a/EX_rs2 [4], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b24/and_b0_9  (\t/a/aluin/sel1_b24/B9 , \t/a/aluin/o_B1 [24], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b24/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b24/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b24/B2 , \t/a/aluin/sel1_b24/B3 );
  or \t/a/aluin/sel1_b24/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b24/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b24/or_B8_B9_o );
  or \t/a/aluin/sel1_b24/or_B8_B9  (\t/a/aluin/sel1_b24/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b24/B9 );
  or \t/a/aluin/sel1_b24/or_or_or_B0_B1_o_or_  (\t/a/EX_B [24], \t/a/aluin/sel1_b24/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b24/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b25/and_b0_2  (\t/a/aluin/sel1_b25/B2 , \t/a/EX_fun7 [0], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b25/and_b0_3  (\t/a/aluin/sel1_b25/B3 , \t/a/EX_fun7 [0], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b25/and_b0_9  (\t/a/aluin/sel1_b25/B9 , \t/a/aluin/o_B1 [25], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b25/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b25/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b25/B2 , \t/a/aluin/sel1_b25/B3 );
  or \t/a/aluin/sel1_b25/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b25/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b25/or_B8_B9_o );
  or \t/a/aluin/sel1_b25/or_B8_B9  (\t/a/aluin/sel1_b25/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b25/B9 );
  or \t/a/aluin/sel1_b25/or_or_or_B0_B1_o_or_  (\t/a/EX_B [25], \t/a/aluin/sel1_b25/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b25/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b26/and_b0_2  (\t/a/aluin/sel1_b26/B2 , \t/a/EX_fun7 [1], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b26/and_b0_3  (\t/a/aluin/sel1_b26/B3 , \t/a/EX_fun7 [1], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b26/and_b0_9  (\t/a/aluin/sel1_b26/B9 , \t/a/aluin/o_B1 [26], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b26/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b26/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b26/B2 , \t/a/aluin/sel1_b26/B3 );
  or \t/a/aluin/sel1_b26/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b26/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b26/or_B8_B9_o );
  or \t/a/aluin/sel1_b26/or_B8_B9  (\t/a/aluin/sel1_b26/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b26/B9 );
  or \t/a/aluin/sel1_b26/or_or_or_B0_B1_o_or_  (\t/a/EX_B [26], \t/a/aluin/sel1_b26/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b26/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b27/and_b0_2  (\t/a/aluin/sel1_b27/B2 , \t/a/EX_fun7 [2], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b27/and_b0_3  (\t/a/aluin/sel1_b27/B3 , \t/a/EX_fun7 [2], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b27/and_b0_9  (\t/a/aluin/sel1_b27/B9 , \t/a/aluin/o_B1 [27], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b27/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b27/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b27/B2 , \t/a/aluin/sel1_b27/B3 );
  or \t/a/aluin/sel1_b27/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b27/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b27/or_B8_B9_o );
  or \t/a/aluin/sel1_b27/or_B8_B9  (\t/a/aluin/sel1_b27/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b27/B9 );
  or \t/a/aluin/sel1_b27/or_or_or_B0_B1_o_or_  (\t/a/EX_B [27], \t/a/aluin/sel1_b27/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b27/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b28/and_b0_2  (\t/a/aluin/sel1_b28/B2 , \t/a/EX_fun7 [3], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b28/and_b0_3  (\t/a/aluin/sel1_b28/B3 , \t/a/EX_fun7 [3], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b28/and_b0_9  (\t/a/aluin/sel1_b28/B9 , \t/a/aluin/o_B1 [28], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b28/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b28/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b28/B2 , \t/a/aluin/sel1_b28/B3 );
  or \t/a/aluin/sel1_b28/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b28/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b28/or_B8_B9_o );
  or \t/a/aluin/sel1_b28/or_B8_B9  (\t/a/aluin/sel1_b28/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b28/B9 );
  or \t/a/aluin/sel1_b28/or_or_or_B0_B1_o_or_  (\t/a/EX_B [28], \t/a/aluin/sel1_b28/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b28/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b29/and_b0_2  (\t/a/aluin/sel1_b29/B2 , \t/a/EX_fun7 [4], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b29/and_b0_3  (\t/a/aluin/sel1_b29/B3 , \t/a/EX_fun7 [4], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b29/and_b0_9  (\t/a/aluin/sel1_b29/B9 , \t/a/aluin/o_B1 [29], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b29/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b29/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b29/B2 , \t/a/aluin/sel1_b29/B3 );
  or \t/a/aluin/sel1_b29/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b29/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b29/or_B8_B9_o );
  or \t/a/aluin/sel1_b29/or_B8_B9  (\t/a/aluin/sel1_b29/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b29/B9 );
  or \t/a/aluin/sel1_b29/or_or_or_B0_B1_o_or_  (\t/a/EX_B [29], \t/a/aluin/sel1_b29/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b29/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b3/and_b0_6  (\t/a/aluin/sel1_b3/B6 , \t/a/EX_rs2 [3], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b3/and_b0_7  (\t/a/aluin/sel1_b3/B7 , \t/a/EX_rd [3], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b3/and_b0_8  (\t/a/aluin/sel1_b3/B8 , \t/a/EX_rs2 [3], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b3/and_b0_9  (\t/a/aluin/sel1_b3/B9 , \t/a/aluin/o_B1 [3], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b3/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b3/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b3/B7 , \t/a/aluin/sel1_b3/or_B8_B9_o );
  or \t/a/aluin/sel1_b3/or_B8_B9  (\t/a/aluin/sel1_b3/or_B8_B9_o , \t/a/aluin/sel1_b3/B8 , \t/a/aluin/sel1_b3/B9 );
  or \t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b3/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b3/B6 , \t/a/aluin/sel1_b3/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b30/and_b0_2  (\t/a/aluin/sel1_b30/B2 , \t/a/EX_fun7 [5], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b30/and_b0_3  (\t/a/aluin/sel1_b30/B3 , \t/a/EX_fun7 [5], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b30/and_b0_9  (\t/a/aluin/sel1_b30/B9 , \t/a/aluin/o_B1 [30], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b30/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b30/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b30/B2 , \t/a/aluin/sel1_b30/B3 );
  or \t/a/aluin/sel1_b30/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b30/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b30/or_B8_B9_o );
  or \t/a/aluin/sel1_b30/or_B8_B9  (\t/a/aluin/sel1_b30/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b30/B9 );
  or \t/a/aluin/sel1_b30/or_or_or_B0_B1_o_or_  (\t/a/EX_B [30], \t/a/aluin/sel1_b30/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b30/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b31/and_b0_2  (\t/a/aluin/sel1_b31/B2 , \t/a/EX_fun7 [6], \t/a/aluin/n4 );
  and \t/a/aluin/sel1_b31/and_b0_3  (\t/a/aluin/sel1_b31/B3 , \t/a/EX_fun7 [6], \t/a/aluin/n1 );
  and \t/a/aluin/sel1_b31/and_b0_9  (\t/a/aluin/sel1_b31/B9 , \t/a/aluin/o_B1 [31], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b31/or_B2_or_B3_B4_o  (\t/a/aluin/sel1_b31/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b31/B2 , \t/a/aluin/sel1_b31/B3 );
  or \t/a/aluin/sel1_b31/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b31/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b11/B7 , \t/a/aluin/sel1_b31/or_B8_B9_o );
  or \t/a/aluin/sel1_b31/or_B8_B9  (\t/a/aluin/sel1_b31/or_B8_B9_o , \t/a/aluin/sel1_b11/B8 , \t/a/aluin/sel1_b31/B9 );
  or \t/a/aluin/sel1_b31/or_or_or_B0_B1_o_or_  (\t/a/EX_B [31], \t/a/aluin/sel1_b31/or_B2_or_B3_B4_o_o , \t/a/aluin/sel1_b31/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b4/and_b0_6  (\t/a/aluin/sel1_b4/B6 , \t/a/EX_rs2 [4], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b4/and_b0_7  (\t/a/aluin/sel1_b4/B7 , \t/a/EX_rd [4], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b4/and_b0_8  (\t/a/aluin/sel1_b4/B8 , \t/a/EX_rs2 [4], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b4/and_b0_9  (\t/a/aluin/sel1_b4/B9 , \t/a/aluin/o_B1 [4], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b4/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b4/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b4/B7 , \t/a/aluin/sel1_b4/or_B8_B9_o );
  or \t/a/aluin/sel1_b4/or_B8_B9  (\t/a/aluin/sel1_b4/or_B8_B9_o , \t/a/aluin/sel1_b4/B8 , \t/a/aluin/sel1_b4/B9 );
  or \t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b4/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b4/B6 , \t/a/aluin/sel1_b4/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b5/and_b0_6  (\t/a/aluin/sel1_b5/B6 , \t/a/aluin/n9 [0], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b5/and_b0_7  (\t/a/aluin/sel1_b5/B7 , \t/a/EX_fun7 [0], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b5/and_b0_8  (\t/a/aluin/sel1_b5/B8 , \t/a/EX_fun7 [0], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b5/and_b0_9  (\t/a/aluin/sel1_b5/B9 , \t/a/aluin/o_B1 [5], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b5/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b5/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b5/B7 , \t/a/aluin/sel1_b5/or_B8_B9_o );
  or \t/a/aluin/sel1_b5/or_B8_B9  (\t/a/aluin/sel1_b5/or_B8_B9_o , \t/a/aluin/sel1_b5/B8 , \t/a/aluin/sel1_b5/B9 );
  or \t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b5/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b5/B6 , \t/a/aluin/sel1_b5/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b6/and_b0_6  (\t/a/aluin/sel1_b6/B6 , \t/a/aluin/n9 [1], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b6/and_b0_7  (\t/a/aluin/sel1_b6/B7 , \t/a/EX_fun7 [1], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b6/and_b0_8  (\t/a/aluin/sel1_b6/B8 , \t/a/EX_fun7 [1], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b6/and_b0_9  (\t/a/aluin/sel1_b6/B9 , \t/a/aluin/o_B1 [6], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b6/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b6/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b6/B7 , \t/a/aluin/sel1_b6/or_B8_B9_o );
  or \t/a/aluin/sel1_b6/or_B8_B9  (\t/a/aluin/sel1_b6/or_B8_B9_o , \t/a/aluin/sel1_b6/B8 , \t/a/aluin/sel1_b6/B9 );
  or \t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b6/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b6/B6 , \t/a/aluin/sel1_b6/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b7/and_b0_6  (\t/a/aluin/sel1_b7/B6 , \t/a/aluin/n9 [2], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b7/and_b0_7  (\t/a/aluin/sel1_b7/B7 , \t/a/EX_fun7 [2], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b7/and_b0_8  (\t/a/aluin/sel1_b7/B8 , \t/a/EX_fun7 [2], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b7/and_b0_9  (\t/a/aluin/sel1_b7/B9 , \t/a/aluin/o_B1 [7], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b7/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b7/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b7/B7 , \t/a/aluin/sel1_b7/or_B8_B9_o );
  or \t/a/aluin/sel1_b7/or_B8_B9  (\t/a/aluin/sel1_b7/or_B8_B9_o , \t/a/aluin/sel1_b7/B8 , \t/a/aluin/sel1_b7/B9 );
  or \t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b7/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b7/B6 , \t/a/aluin/sel1_b7/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b8/and_b0_6  (\t/a/aluin/sel1_b8/B6 , \t/a/aluin/n9 [3], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b8/and_b0_7  (\t/a/aluin/sel1_b8/B7 , \t/a/EX_fun7 [3], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b8/and_b0_8  (\t/a/aluin/sel1_b8/B8 , \t/a/EX_fun7 [3], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b8/and_b0_9  (\t/a/aluin/sel1_b8/B9 , \t/a/aluin/o_B1 [8], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b8/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b8/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b8/B7 , \t/a/aluin/sel1_b8/or_B8_B9_o );
  or \t/a/aluin/sel1_b8/or_B8_B9  (\t/a/aluin/sel1_b8/or_B8_B9_o , \t/a/aluin/sel1_b8/B8 , \t/a/aluin/sel1_b8/B9 );
  or \t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b8/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b8/B6 , \t/a/aluin/sel1_b8/or_B7_or_B8_B9_o_o );
  and \t/a/aluin/sel1_b9/and_b0_6  (\t/a/aluin/sel1_b9/B6 , \t/a/aluin/n9 [4], \t/a/aluin/n13 );
  and \t/a/aluin/sel1_b9/and_b0_7  (\t/a/aluin/sel1_b9/B7 , \t/a/EX_fun7 [4], \t/a/aluin/n12 );
  and \t/a/aluin/sel1_b9/and_b0_8  (\t/a/aluin/sel1_b9/B8 , \t/a/EX_fun7 [4], \t/a/aluin/n11 );
  and \t/a/aluin/sel1_b9/and_b0_9  (\t/a/aluin/sel1_b9/B9 , \t/a/aluin/o_B1 [9], \t/a/aluin/n10 );
  or \t/a/aluin/sel1_b9/or_B7_or_B8_B9_o  (\t/a/aluin/sel1_b9/or_B7_or_B8_B9_o_o , \t/a/aluin/sel1_b9/B7 , \t/a/aluin/sel1_b9/or_B8_B9_o );
  or \t/a/aluin/sel1_b9/or_B8_B9  (\t/a/aluin/sel1_b9/or_B8_B9_o , \t/a/aluin/sel1_b9/B8 , \t/a/aluin/sel1_b9/B9 );
  or \t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7_  (\t/a/aluin/sel1_b9/or_or_B5_B6_o_or_B7__o , \t/a/aluin/sel1_b9/B6 , \t/a/aluin/sel1_b9/or_B7_or_B8_B9_o_o );
  AL_MUX \t/a/aluin/sel2_b0  (
    .i0(1'b0),
    .i1(\t/a/aluin/operation_R [0]),
    .sel(\t/a/aluin/sel2_b0_sel_o ),
    .o(\t/a/EX_operation [0]));  // alu.v(89)
  or \t/a/aluin/sel2_b0_sel  (\t/a/aluin/sel2_b0_sel_o , \t/a/aluin/n13 , \t/a/aluin/n10 );  // alu.v(89)
  AL_MUX \t/a/aluin/sel2_b1  (
    .i0(1'b0),
    .i1(\t/a/EX_fun3 [1]),
    .sel(\t/a/aluin/sel2_b1_sel_is_1_o ),
    .o(\t/a/EX_operation [1]));
  and \t/a/aluin/sel2_b1_sel_is_1  (\t/a/aluin/sel2_b1_sel_is_1_o , \t/a/aluin/sel2_b0_sel_o , \t/a/aluin/mux4_b1_sel_is_1_o_neg );
  AL_MUX \t/a/aluin/sel2_b2  (
    .i0(1'b0),
    .i1(\t/a/aluin/operation_R [2]),
    .sel(\t/a/aluin/sel2_b0_sel_o ),
    .o(\t/a/EX_operation [2]));  // alu.v(89)
  AL_MUX \t/a/aluin/sel2_b3  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\t/a/aluin/sel2_b3_sel_is_3_o ),
    .o(\t/a/EX_operation [3]));
  and \t/a/aluin/sel2_b3_sel_is_3  (\t/a/aluin/sel2_b3_sel_is_3_o , \t/a/aluin/sel2_b0_sel_o , \t/a/aluin/mux4_b1_sel_is_1_o );
  not \t/a/aluin/u2  (\t/a/aluin/n5 , \t/a/aluin/n0 );  // alu.v(54)
  and \t/a/aluin/u23  (\t/a/aluin/n34 , \t/a/aluin/n32 , \t/a/aluin/n10 );  // alu.v(94)
  and \t/a/aluin/u24  (\t/a/aluin/n36 , \t/a/aluin/n34 , \t/a/aluin/n35 );  // alu.v(94)
  and \t/a/aluin/u27  (\t/a/aluin/n39 , \t/a/aluin/n7 , \t/a/aluin/n35 );  // alu.v(96)
  or \t/a/aluin/u3  (\t/a/aluin/n0 , \t/a/aluin/n15 , \t/a/aluin/n14 );  // alu.v(54)
  or \t/a/aluin/u4  (\t/a/aluin/n8 , \t/a/aluin/n6 , \t/a/aluin/n7 );  // alu.v(64)
  or \t/a/aluin/u5  (\t/a/aluin/n14 , \t/a/aluin/n2 , \t/a/aluin/n1 );  // alu.v(54)
  or \t/a/aluin/u9  (\t/a/aluin/n15 , \t/a/aluin/n4 , \t/a/aluin/n3 );  // alu.v(54)
  add_pu32_pu32_o32 \t/a/condition/add0  (
    .i0({\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 [6],\t/a/ID_fun7 ,\t/a/ID_rs2 }),
    .i1(\t/a/ID_jump_regdat1 ),
    .o({\t/a/condition/n5 [31:1],open_n0}));  // PC.v(291)
  eq_w1 \t/a/condition/eq0  (
    .i0(\t/a/ID_jump_risk_block ),
    .i1(1'b1),
    .o(\t/a/condition/n0 ));  // PC.v(266)
  eq_w7 \t/a/condition/eq1  (
    .i0(\t/a/ID_op ),
    .i1(7'b1100111),
    .o(\t/a/condition/JALR_jump_cs ));  // PC.v(272)
  eq_w7 \t/a/condition/eq2  (
    .i0(\t/a/ID_op ),
    .i1(7'b1100011),
    .o(\t/a/condition/n1 ));  // PC.v(276)
  eq_w32 \t/a/condition/eq3  (
    .i0(\t/a/ID_jump_regdat1 ),
    .i1(\t/a/ID_jump_regdat2 ),
    .o(\t/a/condition/n7 ));  // PC.v(312)
  lt_u32_u32 \t/a/condition/lt0  (
    .ci(1'b0),
    .i0(\t/a/ID_jump_regdat1 ),
    .i1(\t/a/ID_jump_regdat2 ),
    .o(\t/a/condition/n9 ));  // PC.v(314)
  lt_u31_u31 \t/a/condition/lt1  (
    .ci(1'b0),
    .i0(\t/a/ID_jump_regdat1 [30:0]),
    .i1(\t/a/ID_jump_regdat2 [30:0]),
    .o(\t/a/condition/n10 ));  // PC.v(315)
  binary_mux_s1_w1 \t/a/condition/mux0_b1  (
    .i0(\t/a/condition/sel0_b1/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [1]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b10  (
    .i0(\t/a/condition/sel0_b10/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [10]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b11  (
    .i0(\t/a/condition/sel0_b11/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [11]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b12  (
    .i0(\t/a/condition/sel0_b12/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [12]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b13  (
    .i0(\t/a/condition/sel0_b13/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [13]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b14  (
    .i0(\t/a/condition/sel0_b14/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [14]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b15  (
    .i0(\t/a/condition/sel0_b15/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [15]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b16  (
    .i0(\t/a/condition/sel0_b16/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [16]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b17  (
    .i0(\t/a/condition/sel0_b17/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [17]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b18  (
    .i0(\t/a/condition/sel0_b18/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [18]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b19  (
    .i0(\t/a/condition/sel0_b19/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [19]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b2  (
    .i0(\t/a/condition/sel0_b2/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [2]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b20  (
    .i0(\t/a/condition/sel0_b20/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [20]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b21  (
    .i0(\t/a/condition/sel0_b21/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [21]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b22  (
    .i0(\t/a/condition/sel0_b22/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [22]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b23  (
    .i0(\t/a/condition/sel0_b23/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [23]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b24  (
    .i0(\t/a/condition/sel0_b24/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [24]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b25  (
    .i0(\t/a/condition/sel0_b25/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [25]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b26  (
    .i0(\t/a/condition/sel0_b26/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [26]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b27  (
    .i0(\t/a/condition/sel0_b27/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [27]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b28  (
    .i0(\t/a/condition/sel0_b28/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [28]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b29  (
    .i0(\t/a/condition/sel0_b29/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [29]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b3  (
    .i0(\t/a/condition/sel0_b3/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [3]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b30  (
    .i0(\t/a/condition/sel0_b30/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [30]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b31  (
    .i0(\t/a/condition/sel0_b31/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [31]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b4  (
    .i0(\t/a/condition/sel0_b4/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [4]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b5  (
    .i0(\t/a/condition/sel0_b5/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [5]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b6  (
    .i0(\t/a/condition/sel0_b6/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [6]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b7  (
    .i0(\t/a/condition/sel0_b7/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [7]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b8  (
    .i0(\t/a/condition/sel0_b8/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [8]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux0_b9  (
    .i0(\t/a/condition/sel0_b9/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_addr [9]));  // PC.v(285)
  binary_mux_s1_w1 \t/a/condition/mux1_b1  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [1]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [1]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b10  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [10]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [10]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b11  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [11]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [11]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b12  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [12]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [12]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b13  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [13]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [13]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b14  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [14]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [14]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b15  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [15]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [15]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b16  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [16]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [16]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b17  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [17]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [17]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b18  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [18]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [18]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b19  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [19]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [19]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b2  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [2]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [2]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b20  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [20]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [20]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b21  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [21]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [21]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b22  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [22]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [22]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b23  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [23]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [23]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b24  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [24]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [24]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b25  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [25]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [25]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b26  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [26]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [26]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b27  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [27]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [27]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b28  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [28]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [28]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b29  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [29]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [29]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b3  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [3]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [3]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b30  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [30]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [30]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b31  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [31]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [31]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b4  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [4]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [4]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b5  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [5]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [5]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b6  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [6]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [6]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b7  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [7]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [7]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b8  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [8]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [8]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux1_b9  (
    .i0(1'b0),
    .i1(\t/a/condition/n5 [9]),
    .sel(\t/a/condition/JALR_jump_cs ),
    .o(\t/a/condition/JALR_jump_addr [9]));  // PC.v(297)
  binary_mux_s1_w1 \t/a/condition/mux2_b1  (
    .i0(1'b0),
    .i1(\t/a/ID_rd [1]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [1]));  // PC.v(306)
  binary_mux_s1_w1 \t/a/condition/mux2_b10  (
    .i0(1'b0),
    .i1(\t/a/ID_fun7 [5]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [10]));  // PC.v(306)
  binary_mux_s1_w1 \t/a/condition/mux2_b11  (
    .i0(1'b0),
    .i1(\t/a/ID_rd [0]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [11]));  // PC.v(306)
  binary_mux_s1_w1 \t/a/condition/mux2_b12  (
    .i0(1'b0),
    .i1(\t/a/ID_fun7 [6]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [12]));  // PC.v(306)
  binary_mux_s1_w1 \t/a/condition/mux2_b2  (
    .i0(1'b0),
    .i1(\t/a/ID_rd [2]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [2]));  // PC.v(306)
  binary_mux_s1_w1 \t/a/condition/mux2_b3  (
    .i0(1'b0),
    .i1(\t/a/ID_rd [3]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [3]));  // PC.v(306)
  binary_mux_s1_w1 \t/a/condition/mux2_b4  (
    .i0(1'b0),
    .i1(\t/a/ID_rd [4]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [4]));  // PC.v(306)
  binary_mux_s1_w1 \t/a/condition/mux2_b5  (
    .i0(1'b0),
    .i1(\t/a/ID_fun7 [0]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [5]));  // PC.v(306)
  binary_mux_s1_w1 \t/a/condition/mux2_b6  (
    .i0(1'b0),
    .i1(\t/a/ID_fun7 [1]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [6]));  // PC.v(306)
  binary_mux_s1_w1 \t/a/condition/mux2_b7  (
    .i0(1'b0),
    .i1(\t/a/ID_fun7 [2]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [7]));  // PC.v(306)
  binary_mux_s1_w1 \t/a/condition/mux2_b8  (
    .i0(1'b0),
    .i1(\t/a/ID_fun7 [3]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [8]));  // PC.v(306)
  binary_mux_s1_w1 \t/a/condition/mux2_b9  (
    .i0(1'b0),
    .i1(\t/a/ID_fun7 [4]),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_addr [9]));  // PC.v(306)
  binary_mux_s3_w1 \t/a/condition/mux3  (
    .i0(\t/a/condition/n7 ),
    .i1(\t/a/condition/n8 ),
    .i2(1'b0),
    .i3(1'b0),
    .i4(\t/a/condition/n9 ),
    .i5(\t/a/condition/n11 ),
    .i6(\t/a/condition/n10 ),
    .i7(\t/a/condition/n12 ),
    .sel(\t/a/ID_fun3 ),
    .o(\t/a/condition/n13 ));  // PC.v(319)
  ne_w32 \t/a/condition/neq0  (
    .i0(\t/a/ID_jump_regdat1 ),
    .i1(\t/a/ID_jump_regdat2 ),
    .o(\t/a/condition/n8 ));  // PC.v(313)
  and \t/a/condition/sel0_b1/and_b0_1  (\t/a/condition/sel0_b1/B1 , \t/a/condition/SB_jump_addr [1], \t/a/condition/n1 );
  and \t/a/condition/sel0_b1/and_b0_2  (\t/a/condition/sel0_b1/B2 , \t/a/condition/JALR_jump_addr [1], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b1/or_B1_B2  (\t/a/condition/sel0_b1/or_B1_B2_o , \t/a/condition/sel0_b1/B1 , \t/a/condition/sel0_b1/B2 );
  and \t/a/condition/sel0_b10/and_b0_1  (\t/a/condition/sel0_b10/B1 , \t/a/condition/SB_jump_addr [10], \t/a/condition/n1 );
  and \t/a/condition/sel0_b10/and_b0_2  (\t/a/condition/sel0_b10/B2 , \t/a/condition/JALR_jump_addr [10], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b10/or_B1_B2  (\t/a/condition/sel0_b10/or_B1_B2_o , \t/a/condition/sel0_b10/B1 , \t/a/condition/sel0_b10/B2 );
  and \t/a/condition/sel0_b11/and_b0_1  (\t/a/condition/sel0_b11/B1 , \t/a/condition/SB_jump_addr [11], \t/a/condition/n1 );
  and \t/a/condition/sel0_b11/and_b0_2  (\t/a/condition/sel0_b11/B2 , \t/a/condition/JALR_jump_addr [11], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b11/or_B1_B2  (\t/a/condition/sel0_b11/or_B1_B2_o , \t/a/condition/sel0_b11/B1 , \t/a/condition/sel0_b11/B2 );
  and \t/a/condition/sel0_b12/and_b0_1  (\t/a/condition/sel0_b12/B1 , \t/a/condition/SB_jump_addr [12], \t/a/condition/n1 );
  and \t/a/condition/sel0_b12/and_b0_2  (\t/a/condition/sel0_b12/B2 , \t/a/condition/JALR_jump_addr [12], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b12/or_B1_B2  (\t/a/condition/sel0_b12/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b12/B2 );
  and \t/a/condition/sel0_b13/and_b0_2  (\t/a/condition/sel0_b13/B2 , \t/a/condition/JALR_jump_addr [13], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b13/or_B1_B2  (\t/a/condition/sel0_b13/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b13/B2 );
  and \t/a/condition/sel0_b14/and_b0_2  (\t/a/condition/sel0_b14/B2 , \t/a/condition/JALR_jump_addr [14], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b14/or_B1_B2  (\t/a/condition/sel0_b14/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b14/B2 );
  and \t/a/condition/sel0_b15/and_b0_2  (\t/a/condition/sel0_b15/B2 , \t/a/condition/JALR_jump_addr [15], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b15/or_B1_B2  (\t/a/condition/sel0_b15/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b15/B2 );
  and \t/a/condition/sel0_b16/and_b0_2  (\t/a/condition/sel0_b16/B2 , \t/a/condition/JALR_jump_addr [16], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b16/or_B1_B2  (\t/a/condition/sel0_b16/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b16/B2 );
  and \t/a/condition/sel0_b17/and_b0_2  (\t/a/condition/sel0_b17/B2 , \t/a/condition/JALR_jump_addr [17], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b17/or_B1_B2  (\t/a/condition/sel0_b17/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b17/B2 );
  and \t/a/condition/sel0_b18/and_b0_2  (\t/a/condition/sel0_b18/B2 , \t/a/condition/JALR_jump_addr [18], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b18/or_B1_B2  (\t/a/condition/sel0_b18/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b18/B2 );
  and \t/a/condition/sel0_b19/and_b0_2  (\t/a/condition/sel0_b19/B2 , \t/a/condition/JALR_jump_addr [19], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b19/or_B1_B2  (\t/a/condition/sel0_b19/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b19/B2 );
  and \t/a/condition/sel0_b2/and_b0_1  (\t/a/condition/sel0_b2/B1 , \t/a/condition/SB_jump_addr [2], \t/a/condition/n1 );
  and \t/a/condition/sel0_b2/and_b0_2  (\t/a/condition/sel0_b2/B2 , \t/a/condition/JALR_jump_addr [2], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b2/or_B1_B2  (\t/a/condition/sel0_b2/or_B1_B2_o , \t/a/condition/sel0_b2/B1 , \t/a/condition/sel0_b2/B2 );
  and \t/a/condition/sel0_b20/and_b0_2  (\t/a/condition/sel0_b20/B2 , \t/a/condition/JALR_jump_addr [20], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b20/or_B1_B2  (\t/a/condition/sel0_b20/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b20/B2 );
  and \t/a/condition/sel0_b21/and_b0_2  (\t/a/condition/sel0_b21/B2 , \t/a/condition/JALR_jump_addr [21], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b21/or_B1_B2  (\t/a/condition/sel0_b21/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b21/B2 );
  and \t/a/condition/sel0_b22/and_b0_2  (\t/a/condition/sel0_b22/B2 , \t/a/condition/JALR_jump_addr [22], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b22/or_B1_B2  (\t/a/condition/sel0_b22/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b22/B2 );
  and \t/a/condition/sel0_b23/and_b0_2  (\t/a/condition/sel0_b23/B2 , \t/a/condition/JALR_jump_addr [23], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b23/or_B1_B2  (\t/a/condition/sel0_b23/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b23/B2 );
  and \t/a/condition/sel0_b24/and_b0_2  (\t/a/condition/sel0_b24/B2 , \t/a/condition/JALR_jump_addr [24], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b24/or_B1_B2  (\t/a/condition/sel0_b24/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b24/B2 );
  and \t/a/condition/sel0_b25/and_b0_2  (\t/a/condition/sel0_b25/B2 , \t/a/condition/JALR_jump_addr [25], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b25/or_B1_B2  (\t/a/condition/sel0_b25/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b25/B2 );
  and \t/a/condition/sel0_b26/and_b0_2  (\t/a/condition/sel0_b26/B2 , \t/a/condition/JALR_jump_addr [26], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b26/or_B1_B2  (\t/a/condition/sel0_b26/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b26/B2 );
  and \t/a/condition/sel0_b27/and_b0_2  (\t/a/condition/sel0_b27/B2 , \t/a/condition/JALR_jump_addr [27], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b27/or_B1_B2  (\t/a/condition/sel0_b27/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b27/B2 );
  and \t/a/condition/sel0_b28/and_b0_2  (\t/a/condition/sel0_b28/B2 , \t/a/condition/JALR_jump_addr [28], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b28/or_B1_B2  (\t/a/condition/sel0_b28/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b28/B2 );
  and \t/a/condition/sel0_b29/and_b0_2  (\t/a/condition/sel0_b29/B2 , \t/a/condition/JALR_jump_addr [29], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b29/or_B1_B2  (\t/a/condition/sel0_b29/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b29/B2 );
  and \t/a/condition/sel0_b3/and_b0_1  (\t/a/condition/sel0_b3/B1 , \t/a/condition/SB_jump_addr [3], \t/a/condition/n1 );
  and \t/a/condition/sel0_b3/and_b0_2  (\t/a/condition/sel0_b3/B2 , \t/a/condition/JALR_jump_addr [3], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b3/or_B1_B2  (\t/a/condition/sel0_b3/or_B1_B2_o , \t/a/condition/sel0_b3/B1 , \t/a/condition/sel0_b3/B2 );
  and \t/a/condition/sel0_b30/and_b0_2  (\t/a/condition/sel0_b30/B2 , \t/a/condition/JALR_jump_addr [30], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b30/or_B1_B2  (\t/a/condition/sel0_b30/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b30/B2 );
  and \t/a/condition/sel0_b31/and_b0_2  (\t/a/condition/sel0_b31/B2 , \t/a/condition/JALR_jump_addr [31], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b31/or_B1_B2  (\t/a/condition/sel0_b31/or_B1_B2_o , \t/a/condition/sel0_b12/B1 , \t/a/condition/sel0_b31/B2 );
  and \t/a/condition/sel0_b4/and_b0_1  (\t/a/condition/sel0_b4/B1 , \t/a/condition/SB_jump_addr [4], \t/a/condition/n1 );
  and \t/a/condition/sel0_b4/and_b0_2  (\t/a/condition/sel0_b4/B2 , \t/a/condition/JALR_jump_addr [4], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b4/or_B1_B2  (\t/a/condition/sel0_b4/or_B1_B2_o , \t/a/condition/sel0_b4/B1 , \t/a/condition/sel0_b4/B2 );
  and \t/a/condition/sel0_b5/and_b0_1  (\t/a/condition/sel0_b5/B1 , \t/a/condition/SB_jump_addr [5], \t/a/condition/n1 );
  and \t/a/condition/sel0_b5/and_b0_2  (\t/a/condition/sel0_b5/B2 , \t/a/condition/JALR_jump_addr [5], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b5/or_B1_B2  (\t/a/condition/sel0_b5/or_B1_B2_o , \t/a/condition/sel0_b5/B1 , \t/a/condition/sel0_b5/B2 );
  and \t/a/condition/sel0_b6/and_b0_1  (\t/a/condition/sel0_b6/B1 , \t/a/condition/SB_jump_addr [6], \t/a/condition/n1 );
  and \t/a/condition/sel0_b6/and_b0_2  (\t/a/condition/sel0_b6/B2 , \t/a/condition/JALR_jump_addr [6], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b6/or_B1_B2  (\t/a/condition/sel0_b6/or_B1_B2_o , \t/a/condition/sel0_b6/B1 , \t/a/condition/sel0_b6/B2 );
  and \t/a/condition/sel0_b7/and_b0_1  (\t/a/condition/sel0_b7/B1 , \t/a/condition/SB_jump_addr [7], \t/a/condition/n1 );
  and \t/a/condition/sel0_b7/and_b0_2  (\t/a/condition/sel0_b7/B2 , \t/a/condition/JALR_jump_addr [7], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b7/or_B1_B2  (\t/a/condition/sel0_b7/or_B1_B2_o , \t/a/condition/sel0_b7/B1 , \t/a/condition/sel0_b7/B2 );
  and \t/a/condition/sel0_b8/and_b0_1  (\t/a/condition/sel0_b8/B1 , \t/a/condition/SB_jump_addr [8], \t/a/condition/n1 );
  and \t/a/condition/sel0_b8/and_b0_2  (\t/a/condition/sel0_b8/B2 , \t/a/condition/JALR_jump_addr [8], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b8/or_B1_B2  (\t/a/condition/sel0_b8/or_B1_B2_o , \t/a/condition/sel0_b8/B1 , \t/a/condition/sel0_b8/B2 );
  and \t/a/condition/sel0_b9/and_b0_1  (\t/a/condition/sel0_b9/B1 , \t/a/condition/SB_jump_addr [9], \t/a/condition/n1 );
  and \t/a/condition/sel0_b9/and_b0_2  (\t/a/condition/sel0_b9/B2 , \t/a/condition/JALR_jump_addr [9], \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel0_b9/or_B1_B2  (\t/a/condition/sel0_b9/or_B1_B2_o , \t/a/condition/sel0_b9/B1 , \t/a/condition/sel0_b9/B2 );
  and \t/a/condition/sel1/and_b0_1  (\t/a/condition/sel1/B1 , \t/a/condition/SB_jump_cs , \t/a/condition/n1 );
  and \t/a/condition/sel1/and_b0_2  (\t/a/condition/sel1/B2 , \t/a/condition/JALR_jump_cs , \t/a/condition/JALR_jump_cs );
  or \t/a/condition/sel1/or_B1_B2  (\t/a/condition/sel1/or_B1_B2_o , \t/a/condition/sel1/B1 , \t/a/condition/sel1/B2 );
  AL_MUX \t/a/condition/u2  (
    .i0(\t/a/condition/sel1/or_B1_B2_o ),
    .i1(1'b0),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/ID_jump_cs ));  // PC.v(285)
  not \t/a/condition/u5  (\t/a/condition/n11 , \t/a/condition/n9 );  // PC.v(316)
  not \t/a/condition/u6  (\t/a/condition/n12 , \t/a/condition/n10 );  // PC.v(317)
  AL_MUX \t/a/condition/u7  (
    .i0(1'b0),
    .i1(\t/a/condition/n13 ),
    .sel(\t/a/condition/n1 ),
    .o(\t/a/condition/SB_jump_cs ));  // PC.v(320)
  eq_w7 \t/a/eq0  (
    .i0(\t/a/ID_op ),
    .i1(7'b0000011),
    .o(\t/a/n0 ));  // cpu.v(178)
  eq_w5 \t/a/eq1  (
    .i0(\t/a/ID_rd ),
    .i1(\t/instruction [19:15]),
    .o(\t/a/n3 ));  // cpu.v(180)
  eq_w3 \t/a/eq10  (
    .i0(\t/a/MEM_fun3 ),
    .i1(3'b001),
    .o(\t/a/n36 ));  // cpu.v(298)
  eq_w3 \t/a/eq11  (
    .i0(\t/a/MEM_fun3 ),
    .i1(3'b010),
    .o(\t/a/n37 ));  // cpu.v(299)
  eq_w5 \t/a/eq2  (
    .i0(\t/a/ID_rd ),
    .i1(\t/instruction [24:20]),
    .o(\t/a/n4 ));  // cpu.v(181)
  eq_w5 \t/a/eq3  (
    .i0(\t/a/MEM_rd ),
    .i1(\t/a/EX_rs1 ),
    .o(\t/a/n9 ));  // cpu.v(239)
  eq_w5 \t/a/eq4  (
    .i0(\t/a/WB_rd ),
    .i1(\t/a/EX_rs1 ),
    .o(\t/a/n20 ));  // cpu.v(246)
  eq_w5 \t/a/eq5  (
    .i0(\t/a/MEM_rd ),
    .i1(\t/a/EX_rs2 ),
    .o(\t/a/n24 ));  // cpu.v(256)
  eq_w5 \t/a/eq6  (
    .i0(\t/a/WB_rd ),
    .i1(\t/a/EX_rs2 ),
    .o(\t/a/n28 ));  // cpu.v(263)
  eq_w7 \t/a/eq7  (
    .i0(\t/a/MEM_op ),
    .i1(7'b0000011),
    .o(\t/memread_cs ));  // cpu.v(287)
  eq_w7 \t/a/eq8  (
    .i0(\t/a/MEM_op ),
    .i1(7'b0100011),
    .o(memwrite_cs));  // cpu.v(287)
  eq_w3 \t/a/eq9  (
    .i0(\t/a/MEM_fun3 ),
    .i1(3'b000),
    .o(\t/a/n35 ));  // cpu.v(297)
  reg_ar_as_w1 \t/a/ex_mem/reg0_b0  (
    .clk(clock),
    .d(\t/a/EX_rd [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_rd [0]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg0_b1  (
    .clk(clock),
    .d(\t/a/EX_rd [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_rd [1]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg0_b2  (
    .clk(clock),
    .d(\t/a/EX_rd [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_rd [2]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg0_b3  (
    .clk(clock),
    .d(\t/a/EX_rd [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_rd [3]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg0_b4  (
    .clk(clock),
    .d(\t/a/EX_rd [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_rd [4]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b0  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [0]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b1  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [1]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b10  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [10]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [10]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b11  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [11]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [11]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b12  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [12]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [12]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b13  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [13]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [13]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b14  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [14]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [14]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b15  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [15]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [15]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b16  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [16]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [16]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b17  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [17]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [17]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b18  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [18]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [18]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b19  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [19]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [19]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b2  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [2]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b20  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [20]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [20]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b21  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [21]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [21]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b22  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [22]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [22]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b23  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [23]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [23]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b24  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [24]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [24]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b25  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [25]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [25]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b26  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [26]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [26]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b27  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [27]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [27]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b28  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [28]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [28]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b29  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [29]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [29]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b3  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [3]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b30  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [30]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [30]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b31  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [31]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [31]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b4  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [4]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b5  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [5]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b6  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [6]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b7  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [7]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [7]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b8  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [8]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [8]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg1_b9  (
    .clk(clock),
    .d(\t/a/EX_regdat2 [9]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_regdat2 [9]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg2_b0  (
    .clk(clock),
    .d(\t/a/EX_op [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_op [0]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg2_b1  (
    .clk(clock),
    .d(\t/a/EX_op [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_op [1]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg2_b2  (
    .clk(clock),
    .d(\t/a/EX_op [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_op [2]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg2_b3  (
    .clk(clock),
    .d(\t/a/EX_op [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_op [3]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg2_b4  (
    .clk(clock),
    .d(\t/a/EX_op [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_op [4]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg2_b5  (
    .clk(clock),
    .d(\t/a/EX_op [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_op [5]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg2_b6  (
    .clk(clock),
    .d(\t/a/EX_op [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_op [6]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg3_b0  (
    .clk(clock),
    .d(\t/a/EX_fun3 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_fun3 [0]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg3_b1  (
    .clk(clock),
    .d(\t/a/EX_fun3 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_fun3 [1]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg3_b2  (
    .clk(clock),
    .d(\t/a/EX_fun3 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_fun3 [2]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b0  (
    .clk(clock),
    .d(\t/a/aludat [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [0]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b1  (
    .clk(clock),
    .d(\t/a/aludat [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [1]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b10  (
    .clk(clock),
    .d(\t/a/aludat [10]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [10]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b11  (
    .clk(clock),
    .d(\t/a/aludat [11]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [11]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b12  (
    .clk(clock),
    .d(\t/a/aludat [12]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [12]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b13  (
    .clk(clock),
    .d(\t/a/aludat [13]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [13]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b14  (
    .clk(clock),
    .d(\t/a/aludat [14]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [14]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b15  (
    .clk(clock),
    .d(\t/a/aludat [15]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [15]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b16  (
    .clk(clock),
    .d(\t/a/aludat [16]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [16]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b17  (
    .clk(clock),
    .d(\t/a/aludat [17]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [17]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b18  (
    .clk(clock),
    .d(\t/a/aludat [18]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [18]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b19  (
    .clk(clock),
    .d(\t/a/aludat [19]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [19]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b2  (
    .clk(clock),
    .d(\t/a/aludat [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [2]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b20  (
    .clk(clock),
    .d(\t/a/aludat [20]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [20]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b21  (
    .clk(clock),
    .d(\t/a/aludat [21]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [21]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b22  (
    .clk(clock),
    .d(\t/a/aludat [22]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [22]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b23  (
    .clk(clock),
    .d(\t/a/aludat [23]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [23]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b24  (
    .clk(clock),
    .d(\t/a/aludat [24]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [24]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b25  (
    .clk(clock),
    .d(\t/a/aludat [25]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [25]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b26  (
    .clk(clock),
    .d(\t/a/aludat [26]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [26]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b27  (
    .clk(clock),
    .d(\t/a/aludat [27]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [27]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b28  (
    .clk(clock),
    .d(\t/a/aludat [28]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [28]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b29  (
    .clk(clock),
    .d(\t/a/aludat [29]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [29]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b3  (
    .clk(clock),
    .d(\t/a/aludat [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [3]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b30  (
    .clk(clock),
    .d(\t/a/aludat [30]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [30]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b31  (
    .clk(clock),
    .d(\t/a/aludat [31]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [31]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b4  (
    .clk(clock),
    .d(\t/a/aludat [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [4]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b5  (
    .clk(clock),
    .d(\t/a/aludat [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [5]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b6  (
    .clk(clock),
    .d(\t/a/aludat [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [6]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b7  (
    .clk(clock),
    .d(\t/a/aludat [7]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [7]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b8  (
    .clk(clock),
    .d(\t/a/aludat [8]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [8]));  // flow_line_reg.v(191)
  reg_ar_as_w1 \t/a/ex_mem/reg4_b9  (
    .clk(clock),
    .d(\t/a/aludat [9]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/MEM_aludat [9]));  // flow_line_reg.v(191)
  not \t/a/ex_mem/u10  (\t/a/ex_mem/n0 , rst);  // flow_line_reg.v(176)
  reg_ar_as_w1 \t/a/id_ex/reg0_b0  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [0]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b1  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [1]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b10  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [10]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [10]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b11  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [11]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [11]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b12  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [12]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [12]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b13  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [13]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [13]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b14  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [14]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [14]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b15  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [15]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [15]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b16  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [16]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [16]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b17  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [17]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [17]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b18  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [18]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [18]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b19  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [19]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [19]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b2  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [2]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b20  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [20]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [20]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b21  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [21]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [21]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b22  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [22]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [22]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b23  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [23]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [23]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b24  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [24]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [24]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b25  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [25]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [25]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b26  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [26]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [26]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b27  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [27]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [27]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b28  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [28]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [28]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b29  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [29]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [29]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b3  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [3]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b30  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [30]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [30]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b31  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [31]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [31]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b4  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [4]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b5  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [5]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b6  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [6]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b7  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [7]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [7]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b8  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [8]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [8]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg0_b9  (
    .clk(clock),
    .d(\t/a/ID_read_dat2 [9]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat2 [9]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg1_b0  (
    .clk(clock),
    .d(\t/a/ID_fun3 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_fun3 [0]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg1_b1  (
    .clk(clock),
    .d(\t/a/ID_fun3 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_fun3 [1]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg1_b2  (
    .clk(clock),
    .d(\t/a/ID_fun3 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_fun3 [2]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg2_b0  (
    .clk(clock),
    .d(\t/a/ID_fun7 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_fun7 [0]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg2_b1  (
    .clk(clock),
    .d(\t/a/ID_fun7 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_fun7 [1]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg2_b2  (
    .clk(clock),
    .d(\t/a/ID_fun7 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_fun7 [2]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg2_b3  (
    .clk(clock),
    .d(\t/a/ID_fun7 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_fun7 [3]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg2_b4  (
    .clk(clock),
    .d(\t/a/ID_fun7 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_fun7 [4]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg2_b5  (
    .clk(clock),
    .d(\t/a/ID_fun7 [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_fun7 [5]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg2_b6  (
    .clk(clock),
    .d(\t/a/ID_fun7 [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_fun7 [6]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg3_b0  (
    .clk(clock),
    .d(\t/a/ID_rs2 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rs2 [0]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg3_b1  (
    .clk(clock),
    .d(\t/a/ID_rs2 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rs2 [1]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg3_b2  (
    .clk(clock),
    .d(\t/a/ID_rs2 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rs2 [2]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg3_b3  (
    .clk(clock),
    .d(\t/a/ID_rs2 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rs2 [3]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg3_b4  (
    .clk(clock),
    .d(\t/a/ID_rs2 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rs2 [4]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg4_b0  (
    .clk(clock),
    .d(\t/a/ID_rs1 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rs1 [0]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg4_b1  (
    .clk(clock),
    .d(\t/a/ID_rs1 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rs1 [1]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg4_b2  (
    .clk(clock),
    .d(\t/a/ID_rs1 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rs1 [2]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg4_b3  (
    .clk(clock),
    .d(\t/a/ID_rs1 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rs1 [3]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg4_b4  (
    .clk(clock),
    .d(\t/a/ID_rs1 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rs1 [4]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg5_b0  (
    .clk(clock),
    .d(\t/a/ID_rd [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rd [0]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg5_b1  (
    .clk(clock),
    .d(\t/a/ID_rd [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rd [1]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg5_b2  (
    .clk(clock),
    .d(\t/a/ID_rd [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rd [2]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg5_b3  (
    .clk(clock),
    .d(\t/a/ID_rd [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rd [3]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg5_b4  (
    .clk(clock),
    .d(\t/a/ID_rd [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_rd [4]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg6_b0  (
    .clk(clock),
    .d(\t/a/ID_op [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_op [0]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg6_b1  (
    .clk(clock),
    .d(\t/a/ID_op [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_op [1]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg6_b2  (
    .clk(clock),
    .d(\t/a/ID_op [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_op [2]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg6_b3  (
    .clk(clock),
    .d(\t/a/ID_op [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_op [3]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg6_b4  (
    .clk(clock),
    .d(\t/a/ID_op [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_op [4]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg6_b5  (
    .clk(clock),
    .d(\t/a/ID_op [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_op [5]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg6_b6  (
    .clk(clock),
    .d(\t/a/ID_op [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_op [6]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b0  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [0]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b1  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [1]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b10  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [10]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [10]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b11  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [11]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [11]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b12  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [12]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [12]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b13  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [13]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [13]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b14  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [14]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [14]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b15  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [15]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [15]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b16  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [16]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [16]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b17  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [17]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [17]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b18  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [18]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [18]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b19  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [19]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [19]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b2  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [2]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b20  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [20]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [20]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b21  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [21]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [21]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b22  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [22]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [22]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b23  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [23]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [23]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b24  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [24]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [24]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b25  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [25]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [25]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b26  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [26]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [26]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b27  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [27]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [27]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b28  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [28]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [28]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b29  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [29]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [29]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b3  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [3]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b30  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [30]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [30]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b31  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [31]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [31]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b4  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [4]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b5  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [5]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b6  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [6]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b7  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [7]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [7]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b8  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [8]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [8]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg7_b9  (
    .clk(clock),
    .d(\t/a/ID_memstraddr [9]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_memstraddr [9]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b0  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [0]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b1  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [1]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b10  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [10]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [10]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b11  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [11]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [11]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b12  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [12]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [12]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b13  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [13]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [13]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b14  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [14]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [14]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b15  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [15]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [15]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b16  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [16]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [16]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b17  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [17]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [17]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b18  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [18]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [18]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b19  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [19]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [19]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b2  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [2]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b20  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [20]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [20]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b21  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [21]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [21]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b22  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [22]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [22]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b23  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [23]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [23]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b24  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [24]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [24]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b25  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [25]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [25]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b26  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [26]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [26]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b27  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [27]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [27]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b28  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [28]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [28]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b29  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [29]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [29]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b3  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [3]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b30  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [30]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [30]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b31  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [31]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [31]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b4  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [4]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b5  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [5]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b6  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [6]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b7  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [7]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [7]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b8  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [8]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [8]));  // flow_line_reg.v(139)
  reg_ar_as_w1 \t/a/id_ex/reg8_b9  (
    .clk(clock),
    .d(\t/a/ID_read_dat1 [9]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/EX_regdat1 [9]));  // flow_line_reg.v(139)
  eq_w1 \t/a/if_id/eq0  (
    .i0(\t/instrnop ),
    .i1(1'b1),
    .o(\t/a/if_id/n1 ));  // flow_line_reg.v(51)
  eq_w1 \t/a/if_id/eq1  (
    .i0(\t/bus_block ),
    .i1(1'b1),
    .o(\t/a/if_id/n2 ));  // flow_line_reg.v(52)
  eq_w1 \t/a/if_id/eq2  (
    .i0(\t/a/ID_LW_block ),
    .i1(1'b1),
    .o(\t/a/if_id/n4 ));  // flow_line_reg.v(53)
  eq_w1 \t/a/if_id/eq3  (
    .i0(\t/a/ID_jump_cs ),
    .i1(1'b1),
    .o(\t/a/if_id/n6 ));  // flow_line_reg.v(54)
  binary_mux_s1_w1 \t/a/if_id/mux0_b0  (
    .i0(\t/instruction [0]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n10 [0]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux0_b1  (
    .i0(\t/instruction [1]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n10 [1]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux0_b2  (
    .i0(\t/instruction [2]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n10 [2]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux0_b3  (
    .i0(\t/instruction [3]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n10 [3]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux0_b4  (
    .i0(\t/instruction [4]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n10 [4]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux0_b5  (
    .i0(\t/instruction [5]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n10 [5]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux0_b6  (
    .i0(\t/instruction [6]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n10 [6]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux1_b0  (
    .i0(\t/instruction [12]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n11 [0]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux1_b1  (
    .i0(\t/instruction [13]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n11 [1]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux1_b2  (
    .i0(\t/instruction [14]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n11 [2]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux2_b0  (
    .i0(\t/instruction [25]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n12 [0]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux2_b1  (
    .i0(\t/instruction [26]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n12 [1]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux2_b2  (
    .i0(\t/instruction [27]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n12 [2]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux2_b3  (
    .i0(\t/instruction [28]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n12 [3]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux2_b4  (
    .i0(\t/instruction [29]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n12 [4]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux2_b5  (
    .i0(\t/instruction [30]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n12 [5]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux2_b6  (
    .i0(\t/instruction [31]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n12 [6]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux3_b0  (
    .i0(\t/instruction [7]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n13 [0]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux3_b1  (
    .i0(\t/instruction [8]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n13 [1]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux3_b2  (
    .i0(\t/instruction [9]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n13 [2]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux3_b3  (
    .i0(\t/instruction [10]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n13 [3]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux3_b4  (
    .i0(\t/instruction [11]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n13 [4]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux4_b0  (
    .i0(\t/instruction [15]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n14 [0]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux4_b1  (
    .i0(\t/instruction [16]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n14 [1]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux4_b2  (
    .i0(\t/instruction [17]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n14 [2]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux4_b3  (
    .i0(\t/instruction [18]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n14 [3]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux4_b4  (
    .i0(\t/instruction [19]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n14 [4]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux5_b0  (
    .i0(\t/instruction [20]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n15 [0]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux5_b1  (
    .i0(\t/instruction [21]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n15 [1]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux5_b2  (
    .i0(\t/instruction [22]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n15 [2]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux5_b3  (
    .i0(\t/instruction [23]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n15 [3]));  // flow_line_reg.v(71)
  binary_mux_s1_w1 \t/a/if_id/mux5_b4  (
    .i0(\t/instruction [24]),
    .i1(1'b0),
    .sel(\t/a/if_id/n9 ),
    .o(\t/a/if_id/n15 [4]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg0_b0  (
    .clk(clock),
    .d(\t/a/if_id/n11 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_fun3 [0]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg0_b1  (
    .clk(clock),
    .d(\t/a/if_id/n11 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_fun3 [1]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg0_b2  (
    .clk(clock),
    .d(\t/a/if_id/n11 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_fun3 [2]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg1_b0  (
    .clk(clock),
    .d(\t/a/if_id/n12 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_fun7 [0]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg1_b1  (
    .clk(clock),
    .d(\t/a/if_id/n12 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_fun7 [1]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg1_b2  (
    .clk(clock),
    .d(\t/a/if_id/n12 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_fun7 [2]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg1_b3  (
    .clk(clock),
    .d(\t/a/if_id/n12 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_fun7 [3]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg1_b4  (
    .clk(clock),
    .d(\t/a/if_id/n12 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_fun7 [4]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg1_b5  (
    .clk(clock),
    .d(\t/a/if_id/n12 [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_fun7 [5]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg1_b6  (
    .clk(clock),
    .d(\t/a/if_id/n12 [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_fun7 [6]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg2_b0  (
    .clk(clock),
    .d(\t/a/if_id/n13 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rd [0]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg2_b1  (
    .clk(clock),
    .d(\t/a/if_id/n13 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rd [1]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg2_b2  (
    .clk(clock),
    .d(\t/a/if_id/n13 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rd [2]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg2_b3  (
    .clk(clock),
    .d(\t/a/if_id/n13 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rd [3]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg2_b4  (
    .clk(clock),
    .d(\t/a/if_id/n13 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rd [4]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg3_b0  (
    .clk(clock),
    .d(\t/a/if_id/n14 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rs1 [0]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg3_b1  (
    .clk(clock),
    .d(\t/a/if_id/n14 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rs1 [1]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg3_b2  (
    .clk(clock),
    .d(\t/a/if_id/n14 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rs1 [2]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg3_b3  (
    .clk(clock),
    .d(\t/a/if_id/n14 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rs1 [3]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg3_b4  (
    .clk(clock),
    .d(\t/a/if_id/n14 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rs1 [4]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg4_b0  (
    .clk(clock),
    .d(\t/a/if_id/n15 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rs2 [0]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg4_b1  (
    .clk(clock),
    .d(\t/a/if_id/n15 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rs2 [1]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg4_b2  (
    .clk(clock),
    .d(\t/a/if_id/n15 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rs2 [2]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg4_b3  (
    .clk(clock),
    .d(\t/a/if_id/n15 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rs2 [3]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg4_b4  (
    .clk(clock),
    .d(\t/a/if_id/n15 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_rs2 [4]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b0  (
    .clk(clock),
    .d(\t/memstraddress [0]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [0]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b1  (
    .clk(clock),
    .d(\t/memstraddress [1]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [1]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b10  (
    .clk(clock),
    .d(\t/memstraddress [10]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [10]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b11  (
    .clk(clock),
    .d(\t/memstraddress [11]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [11]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b12  (
    .clk(clock),
    .d(\t/memstraddress [12]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [12]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b13  (
    .clk(clock),
    .d(\t/memstraddress [13]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [13]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b14  (
    .clk(clock),
    .d(\t/memstraddress [14]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [14]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b15  (
    .clk(clock),
    .d(\t/memstraddress [15]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [15]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b16  (
    .clk(clock),
    .d(\t/memstraddress [16]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [16]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b17  (
    .clk(clock),
    .d(\t/memstraddress [17]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [17]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b18  (
    .clk(clock),
    .d(\t/memstraddress [18]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [18]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b19  (
    .clk(clock),
    .d(\t/memstraddress [19]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [19]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b2  (
    .clk(clock),
    .d(\t/memstraddress [2]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [2]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b20  (
    .clk(clock),
    .d(\t/memstraddress [20]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [20]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b21  (
    .clk(clock),
    .d(\t/memstraddress [21]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [21]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b22  (
    .clk(clock),
    .d(\t/memstraddress [22]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [22]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b23  (
    .clk(clock),
    .d(\t/memstraddress [23]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [23]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b24  (
    .clk(clock),
    .d(\t/memstraddress [24]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [24]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b25  (
    .clk(clock),
    .d(\t/memstraddress [25]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [25]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b26  (
    .clk(clock),
    .d(\t/memstraddress [26]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [26]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b27  (
    .clk(clock),
    .d(\t/memstraddress [27]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [27]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b28  (
    .clk(clock),
    .d(\t/memstraddress [28]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [28]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b29  (
    .clk(clock),
    .d(\t/memstraddress [29]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [29]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b3  (
    .clk(clock),
    .d(\t/memstraddress [3]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [3]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b30  (
    .clk(clock),
    .d(\t/memstraddress [30]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [30]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b31  (
    .clk(clock),
    .d(\t/memstraddress [31]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [31]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b4  (
    .clk(clock),
    .d(\t/memstraddress [4]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [4]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b5  (
    .clk(clock),
    .d(\t/memstraddress [5]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [5]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b6  (
    .clk(clock),
    .d(\t/memstraddress [6]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [6]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b7  (
    .clk(clock),
    .d(\t/memstraddress [7]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [7]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b8  (
    .clk(clock),
    .d(\t/memstraddress [8]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [8]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg5_b9  (
    .clk(clock),
    .d(\t/memstraddress [9]),
    .en(~\t/a/if_id/n9 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_memstraddr [9]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg6_b0  (
    .clk(clock),
    .d(\t/a/if_id/n10 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_op [0]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg6_b1  (
    .clk(clock),
    .d(\t/a/if_id/n10 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_op [1]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg6_b2  (
    .clk(clock),
    .d(\t/a/if_id/n10 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_op [2]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg6_b3  (
    .clk(clock),
    .d(\t/a/if_id/n10 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_op [3]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg6_b4  (
    .clk(clock),
    .d(\t/a/if_id/n10 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_op [4]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg6_b5  (
    .clk(clock),
    .d(\t/a/if_id/n10 [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_op [5]));  // flow_line_reg.v(71)
  reg_ar_as_w1 \t/a/if_id/reg6_b6  (
    .clk(clock),
    .d(\t/a/if_id/n10 [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/ID_op [6]));  // flow_line_reg.v(71)
  or \t/a/if_id/u12  (\t/a/if_id/n3 , \t/a/if_id/n1 , \t/a/if_id/n2 );  // flow_line_reg.v(52)
  or \t/a/if_id/u13  (\t/a/if_id/n5 , \t/a/if_id/n3 , \t/a/if_id/n4 );  // flow_line_reg.v(53)
  or \t/a/if_id/u14  (\t/a/if_id/n7 , \t/a/if_id/n5 , \t/a/if_id/n6 );  // flow_line_reg.v(54)
  or \t/a/if_id/u15  (\t/a/if_id/n9 , \t/a/if_id/n7 , \t/a/condition/n0 );  // flow_line_reg.v(55)
  add_pu32_pu32_o32 \t/a/instr/add0  (
    .i0(\t/memstraddress ),
    .i1({\t/a/IF_skip_addr [31:1],1'b0}),
    .o(\t/a/instr/n12 ));  // PC.v(50)
  add_pu32_pu32_o32 \t/a/instr/add1  (
    .i0(\t/memstraddress ),
    .i1({\t/a/ID_jump_addr [31:1],1'b0}),
    .o(\t/a/instr/n14 ));  // PC.v(54)
  add_pu30_pu30_o30 \t/a/instr/add2  (
    .i0(\t/memstraddress [31:2]),
    .i1(30'b000000000000000000000000000001),
    .o(\t/a/instr/n16 ));  // PC.v(58)
  eq_w1 \t/a/instr/eq0  (
    .i0(\t/memread_cs ),
    .i1(1'b1),
    .o(\t/a/instr/n1 ));  // PC.v(35)
  eq_w32 \t/a/instr/eq1  (
    .i0(\t/a/memreaddat ),
    .i1(32'b00000000000000000000000000000000),
    .o(\t/a/instr/n2 ));  // PC.v(35)
  eq_w1 \t/a/instr/eq5  (
    .i0(\t/a/IF_skip_cs ),
    .i1(1'b1),
    .o(\t/a/instr/n11 ));  // PC.v(49)
  reg_ar_as_w1 \t/a/instr/instr_nop_reg  (
    .clk(clock),
    .d(\t/a/instr/n20 ),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/instrnop ));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux0_b0  (
    .i0(\t/memstraddress [0]),
    .i1(\t/a/ID_memstraddr [0]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [0]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b1  (
    .i0(\t/memstraddress [1]),
    .i1(\t/a/ID_memstraddr [1]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [1]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b10  (
    .i0(\t/memstraddress [10]),
    .i1(\t/a/ID_memstraddr [10]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [10]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b11  (
    .i0(\t/memstraddress [11]),
    .i1(\t/a/ID_memstraddr [11]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [11]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b12  (
    .i0(\t/memstraddress [12]),
    .i1(\t/a/ID_memstraddr [12]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [12]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b13  (
    .i0(\t/memstraddress [13]),
    .i1(\t/a/ID_memstraddr [13]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [13]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b14  (
    .i0(\t/memstraddress [14]),
    .i1(\t/a/ID_memstraddr [14]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [14]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b15  (
    .i0(\t/memstraddress [15]),
    .i1(\t/a/ID_memstraddr [15]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [15]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b16  (
    .i0(\t/memstraddress [16]),
    .i1(\t/a/ID_memstraddr [16]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [16]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b17  (
    .i0(\t/memstraddress [17]),
    .i1(\t/a/ID_memstraddr [17]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [17]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b18  (
    .i0(\t/memstraddress [18]),
    .i1(\t/a/ID_memstraddr [18]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [18]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b19  (
    .i0(\t/memstraddress [19]),
    .i1(\t/a/ID_memstraddr [19]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [19]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b2  (
    .i0(\t/memstraddress [2]),
    .i1(\t/a/ID_memstraddr [2]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [2]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b20  (
    .i0(\t/memstraddress [20]),
    .i1(\t/a/ID_memstraddr [20]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [20]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b21  (
    .i0(\t/memstraddress [21]),
    .i1(\t/a/ID_memstraddr [21]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [21]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b22  (
    .i0(\t/memstraddress [22]),
    .i1(\t/a/ID_memstraddr [22]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [22]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b23  (
    .i0(\t/memstraddress [23]),
    .i1(\t/a/ID_memstraddr [23]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [23]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b24  (
    .i0(\t/memstraddress [24]),
    .i1(\t/a/ID_memstraddr [24]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [24]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b25  (
    .i0(\t/memstraddress [25]),
    .i1(\t/a/ID_memstraddr [25]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [25]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b26  (
    .i0(\t/memstraddress [26]),
    .i1(\t/a/ID_memstraddr [26]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [26]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b27  (
    .i0(\t/memstraddress [27]),
    .i1(\t/a/ID_memstraddr [27]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [27]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b28  (
    .i0(\t/memstraddress [28]),
    .i1(\t/a/ID_memstraddr [28]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [28]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b29  (
    .i0(\t/memstraddress [29]),
    .i1(\t/a/ID_memstraddr [29]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [29]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b3  (
    .i0(\t/memstraddress [3]),
    .i1(\t/a/ID_memstraddr [3]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [3]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b30  (
    .i0(\t/memstraddress [30]),
    .i1(\t/a/ID_memstraddr [30]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [30]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b31  (
    .i0(\t/memstraddress [31]),
    .i1(\t/a/ID_memstraddr [31]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [31]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b4  (
    .i0(\t/memstraddress [4]),
    .i1(\t/a/ID_memstraddr [4]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [4]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b5  (
    .i0(\t/memstraddress [5]),
    .i1(\t/a/ID_memstraddr [5]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [5]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b6  (
    .i0(\t/memstraddress [6]),
    .i1(\t/a/ID_memstraddr [6]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [6]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b7  (
    .i0(\t/memstraddress [7]),
    .i1(\t/a/ID_memstraddr [7]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [7]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b8  (
    .i0(\t/memstraddress [8]),
    .i1(\t/a/ID_memstraddr [8]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [8]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux0_b9  (
    .i0(\t/memstraddress [9]),
    .i1(\t/a/ID_memstraddr [9]),
    .sel(\t/a/condition/n0 ),
    .o(\t/a/instr/n10 [9]));  // PC.v(42)
  binary_mux_s1_w1 \t/a/instr/mux1_b0  (
    .i0(\t/memstraddress [0]),
    .i1(\t/a/instr/n15 [0]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [0]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b1  (
    .i0(\t/memstraddress [1]),
    .i1(\t/a/instr/n15 [1]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [1]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b10  (
    .i0(\t/a/instr/n16 [8]),
    .i1(\t/a/instr/n15 [10]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [10]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b11  (
    .i0(\t/a/instr/n16 [9]),
    .i1(\t/a/instr/n15 [11]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [11]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b12  (
    .i0(\t/a/instr/n16 [10]),
    .i1(\t/a/instr/n15 [12]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [12]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b13  (
    .i0(\t/a/instr/n16 [11]),
    .i1(\t/a/instr/n15 [13]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [13]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b14  (
    .i0(\t/a/instr/n16 [12]),
    .i1(\t/a/instr/n15 [14]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [14]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b15  (
    .i0(\t/a/instr/n16 [13]),
    .i1(\t/a/instr/n15 [15]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [15]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b16  (
    .i0(\t/a/instr/n16 [14]),
    .i1(\t/a/instr/n15 [16]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [16]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b17  (
    .i0(\t/a/instr/n16 [15]),
    .i1(\t/a/instr/n15 [17]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [17]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b18  (
    .i0(\t/a/instr/n16 [16]),
    .i1(\t/a/instr/n15 [18]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [18]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b19  (
    .i0(\t/a/instr/n16 [17]),
    .i1(\t/a/instr/n15 [19]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [19]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b2  (
    .i0(\t/a/instr/n16 [0]),
    .i1(\t/a/instr/n15 [2]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [2]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b20  (
    .i0(\t/a/instr/n16 [18]),
    .i1(\t/a/instr/n15 [20]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [20]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b21  (
    .i0(\t/a/instr/n16 [19]),
    .i1(\t/a/instr/n15 [21]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [21]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b22  (
    .i0(\t/a/instr/n16 [20]),
    .i1(\t/a/instr/n15 [22]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [22]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b23  (
    .i0(\t/a/instr/n16 [21]),
    .i1(\t/a/instr/n15 [23]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [23]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b24  (
    .i0(\t/a/instr/n16 [22]),
    .i1(\t/a/instr/n15 [24]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [24]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b25  (
    .i0(\t/a/instr/n16 [23]),
    .i1(\t/a/instr/n15 [25]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [25]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b26  (
    .i0(\t/a/instr/n16 [24]),
    .i1(\t/a/instr/n15 [26]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [26]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b27  (
    .i0(\t/a/instr/n16 [25]),
    .i1(\t/a/instr/n15 [27]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [27]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b28  (
    .i0(\t/a/instr/n16 [26]),
    .i1(\t/a/instr/n15 [28]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [28]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b29  (
    .i0(\t/a/instr/n16 [27]),
    .i1(\t/a/instr/n15 [29]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [29]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b3  (
    .i0(\t/a/instr/n16 [1]),
    .i1(\t/a/instr/n15 [3]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [3]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b30  (
    .i0(\t/a/instr/n16 [28]),
    .i1(\t/a/instr/n15 [30]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [30]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b31  (
    .i0(\t/a/instr/n16 [29]),
    .i1(\t/a/instr/n15 [31]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [31]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b4  (
    .i0(\t/a/instr/n16 [2]),
    .i1(\t/a/instr/n15 [4]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [4]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b5  (
    .i0(\t/a/instr/n16 [3]),
    .i1(\t/a/instr/n15 [5]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [5]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b6  (
    .i0(\t/a/instr/n16 [4]),
    .i1(\t/a/instr/n15 [6]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [6]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b7  (
    .i0(\t/a/instr/n16 [5]),
    .i1(\t/a/instr/n15 [7]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [7]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b8  (
    .i0(\t/a/instr/n16 [6]),
    .i1(\t/a/instr/n15 [8]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [8]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux1_b9  (
    .i0(\t/a/instr/n16 [7]),
    .i1(\t/a/instr/n15 [9]),
    .sel(\t/a/if_id/n6 ),
    .o(\t/a/instr/n17 [9]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b0  (
    .i0(\t/a/instr/n17 [0]),
    .i1(\t/a/instr/n12 [0]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [0]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b1  (
    .i0(\t/a/instr/n17 [1]),
    .i1(\t/a/instr/n12 [1]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [1]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b10  (
    .i0(\t/a/instr/n17 [10]),
    .i1(\t/a/instr/n12 [10]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [10]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b11  (
    .i0(\t/a/instr/n17 [11]),
    .i1(\t/a/instr/n12 [11]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [11]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b12  (
    .i0(\t/a/instr/n17 [12]),
    .i1(\t/a/instr/n12 [12]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [12]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b13  (
    .i0(\t/a/instr/n17 [13]),
    .i1(\t/a/instr/n12 [13]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [13]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b14  (
    .i0(\t/a/instr/n17 [14]),
    .i1(\t/a/instr/n12 [14]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [14]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b15  (
    .i0(\t/a/instr/n17 [15]),
    .i1(\t/a/instr/n12 [15]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [15]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b16  (
    .i0(\t/a/instr/n17 [16]),
    .i1(\t/a/instr/n12 [16]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [16]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b17  (
    .i0(\t/a/instr/n17 [17]),
    .i1(\t/a/instr/n12 [17]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [17]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b18  (
    .i0(\t/a/instr/n17 [18]),
    .i1(\t/a/instr/n12 [18]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [18]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b19  (
    .i0(\t/a/instr/n17 [19]),
    .i1(\t/a/instr/n12 [19]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [19]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b2  (
    .i0(\t/a/instr/n17 [2]),
    .i1(\t/a/instr/n12 [2]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [2]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b20  (
    .i0(\t/a/instr/n17 [20]),
    .i1(\t/a/instr/n12 [20]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [20]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b21  (
    .i0(\t/a/instr/n17 [21]),
    .i1(\t/a/instr/n12 [21]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [21]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b22  (
    .i0(\t/a/instr/n17 [22]),
    .i1(\t/a/instr/n12 [22]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [22]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b23  (
    .i0(\t/a/instr/n17 [23]),
    .i1(\t/a/instr/n12 [23]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [23]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b24  (
    .i0(\t/a/instr/n17 [24]),
    .i1(\t/a/instr/n12 [24]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [24]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b25  (
    .i0(\t/a/instr/n17 [25]),
    .i1(\t/a/instr/n12 [25]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [25]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b26  (
    .i0(\t/a/instr/n17 [26]),
    .i1(\t/a/instr/n12 [26]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [26]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b27  (
    .i0(\t/a/instr/n17 [27]),
    .i1(\t/a/instr/n12 [27]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [27]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b28  (
    .i0(\t/a/instr/n17 [28]),
    .i1(\t/a/instr/n12 [28]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [28]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b29  (
    .i0(\t/a/instr/n17 [29]),
    .i1(\t/a/instr/n12 [29]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [29]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b3  (
    .i0(\t/a/instr/n17 [3]),
    .i1(\t/a/instr/n12 [3]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [3]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b30  (
    .i0(\t/a/instr/n17 [30]),
    .i1(\t/a/instr/n12 [30]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [30]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b31  (
    .i0(\t/a/instr/n17 [31]),
    .i1(\t/a/instr/n12 [31]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [31]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b4  (
    .i0(\t/a/instr/n17 [4]),
    .i1(\t/a/instr/n12 [4]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [4]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b5  (
    .i0(\t/a/instr/n17 [5]),
    .i1(\t/a/instr/n12 [5]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [5]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b6  (
    .i0(\t/a/instr/n17 [6]),
    .i1(\t/a/instr/n12 [6]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [6]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b7  (
    .i0(\t/a/instr/n17 [7]),
    .i1(\t/a/instr/n12 [7]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [7]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b8  (
    .i0(\t/a/instr/n17 [8]),
    .i1(\t/a/instr/n12 [8]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [8]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux2_b9  (
    .i0(\t/a/instr/n17 [9]),
    .i1(\t/a/instr/n12 [9]),
    .sel(\t/a/instr/n11 ),
    .o(\t/a/instr/n18 [9]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b0  (
    .i0(\t/a/instr/n18 [0]),
    .i1(\t/a/instr/n10 [0]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [0]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b1  (
    .i0(\t/a/instr/n18 [1]),
    .i1(\t/a/instr/n10 [1]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [1]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b10  (
    .i0(\t/a/instr/n18 [10]),
    .i1(\t/a/instr/n10 [10]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [10]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b11  (
    .i0(\t/a/instr/n18 [11]),
    .i1(\t/a/instr/n10 [11]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [11]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b12  (
    .i0(\t/a/instr/n18 [12]),
    .i1(\t/a/instr/n10 [12]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [12]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b13  (
    .i0(\t/a/instr/n18 [13]),
    .i1(\t/a/instr/n10 [13]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [13]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b14  (
    .i0(\t/a/instr/n18 [14]),
    .i1(\t/a/instr/n10 [14]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [14]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b15  (
    .i0(\t/a/instr/n18 [15]),
    .i1(\t/a/instr/n10 [15]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [15]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b16  (
    .i0(\t/a/instr/n18 [16]),
    .i1(\t/a/instr/n10 [16]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [16]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b17  (
    .i0(\t/a/instr/n18 [17]),
    .i1(\t/a/instr/n10 [17]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [17]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b18  (
    .i0(\t/a/instr/n18 [18]),
    .i1(\t/a/instr/n10 [18]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [18]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b19  (
    .i0(\t/a/instr/n18 [19]),
    .i1(\t/a/instr/n10 [19]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [19]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b2  (
    .i0(\t/a/instr/n18 [2]),
    .i1(\t/a/instr/n10 [2]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [2]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b20  (
    .i0(\t/a/instr/n18 [20]),
    .i1(\t/a/instr/n10 [20]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [20]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b21  (
    .i0(\t/a/instr/n18 [21]),
    .i1(\t/a/instr/n10 [21]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [21]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b22  (
    .i0(\t/a/instr/n18 [22]),
    .i1(\t/a/instr/n10 [22]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [22]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b23  (
    .i0(\t/a/instr/n18 [23]),
    .i1(\t/a/instr/n10 [23]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [23]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b24  (
    .i0(\t/a/instr/n18 [24]),
    .i1(\t/a/instr/n10 [24]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [24]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b25  (
    .i0(\t/a/instr/n18 [25]),
    .i1(\t/a/instr/n10 [25]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [25]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b26  (
    .i0(\t/a/instr/n18 [26]),
    .i1(\t/a/instr/n10 [26]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [26]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b27  (
    .i0(\t/a/instr/n18 [27]),
    .i1(\t/a/instr/n10 [27]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [27]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b28  (
    .i0(\t/a/instr/n18 [28]),
    .i1(\t/a/instr/n10 [28]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [28]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b29  (
    .i0(\t/a/instr/n18 [29]),
    .i1(\t/a/instr/n10 [29]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [29]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b3  (
    .i0(\t/a/instr/n18 [3]),
    .i1(\t/a/instr/n10 [3]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [3]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b30  (
    .i0(\t/a/instr/n18 [30]),
    .i1(\t/a/instr/n10 [30]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [30]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b31  (
    .i0(\t/a/instr/n18 [31]),
    .i1(\t/a/instr/n10 [31]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [31]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b4  (
    .i0(\t/a/instr/n18 [4]),
    .i1(\t/a/instr/n10 [4]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [4]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b5  (
    .i0(\t/a/instr/n18 [5]),
    .i1(\t/a/instr/n10 [5]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [5]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b6  (
    .i0(\t/a/instr/n18 [6]),
    .i1(\t/a/instr/n10 [6]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [6]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b7  (
    .i0(\t/a/instr/n18 [7]),
    .i1(\t/a/instr/n10 [7]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [7]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b8  (
    .i0(\t/a/instr/n18 [8]),
    .i1(\t/a/instr/n10 [8]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [8]));  // PC.v(60)
  binary_mux_s1_w1 \t/a/instr/mux3_b9  (
    .i0(\t/a/instr/n18 [9]),
    .i1(\t/a/instr/n10 [9]),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n19 [9]));  // PC.v(60)
  not \t/a/instr/n1_inv  (\t/a/instr/n1_neg , \t/a/instr/n1 );
  reg_ar_as_w1 \t/a/instr/reg0_b0  (
    .clk(clock),
    .d(\t/a/instr/n19 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [0]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b1  (
    .clk(clock),
    .d(\t/a/instr/n19 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [1]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b10  (
    .clk(clock),
    .d(\t/a/instr/n19 [10]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [10]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b11  (
    .clk(clock),
    .d(\t/a/instr/n19 [11]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [11]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b12  (
    .clk(clock),
    .d(\t/a/instr/n19 [12]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [12]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b13  (
    .clk(clock),
    .d(\t/a/instr/n19 [13]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [13]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b14  (
    .clk(clock),
    .d(\t/a/instr/n19 [14]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [14]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b15  (
    .clk(clock),
    .d(\t/a/instr/n19 [15]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [15]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b16  (
    .clk(clock),
    .d(\t/a/instr/n19 [16]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [16]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b17  (
    .clk(clock),
    .d(\t/a/instr/n19 [17]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [17]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b18  (
    .clk(clock),
    .d(\t/a/instr/n19 [18]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [18]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b19  (
    .clk(clock),
    .d(\t/a/instr/n19 [19]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [19]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b2  (
    .clk(clock),
    .d(\t/a/instr/n19 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(~rst),
    .q(\t/memstraddress [2]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b20  (
    .clk(clock),
    .d(\t/a/instr/n19 [20]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [20]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b21  (
    .clk(clock),
    .d(\t/a/instr/n19 [21]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [21]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b22  (
    .clk(clock),
    .d(\t/a/instr/n19 [22]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [22]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b23  (
    .clk(clock),
    .d(\t/a/instr/n19 [23]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [23]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b24  (
    .clk(clock),
    .d(\t/a/instr/n19 [24]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [24]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b25  (
    .clk(clock),
    .d(\t/a/instr/n19 [25]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [25]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b26  (
    .clk(clock),
    .d(\t/a/instr/n19 [26]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [26]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b27  (
    .clk(clock),
    .d(\t/a/instr/n19 [27]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [27]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b28  (
    .clk(clock),
    .d(\t/a/instr/n19 [28]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [28]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b29  (
    .clk(clock),
    .d(\t/a/instr/n19 [29]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [29]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b3  (
    .clk(clock),
    .d(\t/a/instr/n19 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [3]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b30  (
    .clk(clock),
    .d(\t/a/instr/n19 [30]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [30]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b31  (
    .clk(clock),
    .d(\t/a/instr/n19 [31]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [31]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b4  (
    .clk(clock),
    .d(\t/a/instr/n19 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [4]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b5  (
    .clk(clock),
    .d(\t/a/instr/n19 [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [5]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b6  (
    .clk(clock),
    .d(\t/a/instr/n19 [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [6]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b7  (
    .clk(clock),
    .d(\t/a/instr/n19 [7]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [7]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b8  (
    .clk(clock),
    .d(\t/a/instr/n19 [8]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [8]));  // PC.v(60)
  reg_ar_as_w1 \t/a/instr/reg0_b9  (
    .clk(clock),
    .d(\t/a/instr/n19 [9]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/memstraddress [9]));  // PC.v(60)
  add_pu32_mu32_o32 \t/a/instr/sub0  (
    .i0(\t/a/instr/n14 ),
    .i1(32'b00000000000000000000000000000100),
    .o(\t/a/instr/n15 ));  // PC.v(54)
  and \t/a/instr/u10  (\t/a/instr/n3 , \t/a/instr/n1 , \t/a/instr/n2 );  // PC.v(35)
  or \t/a/instr/u11  (\t/a/instr/n5 , \t/a/instr/n3 , \t/a/if_id/n4 );  // PC.v(36)
  or \t/a/instr/u12  (\t/a/instr/n7 , \t/a/instr/n5 , \t/a/if_id/n2 );  // PC.v(37)
  or \t/a/instr/u13  (\t/a/instr/n9 , \t/a/instr/n7 , \t/a/condition/n0 );  // PC.v(38)
  AL_MUX \t/a/instr/u18  (
    .i0(1'b0),
    .i1(\t/a/instr/n3 ),
    .sel(\t/a/instr/n9 ),
    .o(\t/a/instr/n20 ));  // PC.v(60)
  eq_w7 \t/a/mem_wb/eq2  (
    .i0(\t/a/MEM_op ),
    .i1(7'b1100011),
    .o(\t/a/mem_wb/n7 ));  // flow_line_reg.v(229)
  eq_w7 \t/a/mem_wb/eq3  (
    .i0(\t/a/MEM_op ),
    .i1(7'b0000000),
    .o(\t/a/mem_wb/n9 ));  // flow_line_reg.v(230)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b0  (
    .i0(\t/a/MEM_aludat [0]),
    .i1(\t/a/memreaddat [0]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [0]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b1  (
    .i0(\t/a/MEM_aludat [1]),
    .i1(\t/a/memreaddat [1]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [1]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b10  (
    .i0(\t/a/MEM_aludat [10]),
    .i1(\t/a/memreaddat [10]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [10]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b11  (
    .i0(\t/a/MEM_aludat [11]),
    .i1(\t/a/memreaddat [11]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [11]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b12  (
    .i0(\t/a/MEM_aludat [12]),
    .i1(\t/a/memreaddat [12]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [12]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b13  (
    .i0(\t/a/MEM_aludat [13]),
    .i1(\t/a/memreaddat [13]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [13]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b14  (
    .i0(\t/a/MEM_aludat [14]),
    .i1(\t/a/memreaddat [14]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [14]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b15  (
    .i0(\t/a/MEM_aludat [15]),
    .i1(\t/a/memreaddat [15]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [15]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b16  (
    .i0(\t/a/MEM_aludat [16]),
    .i1(\t/a/memreaddat [16]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [16]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b17  (
    .i0(\t/a/MEM_aludat [17]),
    .i1(\t/a/memreaddat [17]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [17]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b18  (
    .i0(\t/a/MEM_aludat [18]),
    .i1(\t/a/memreaddat [18]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [18]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b19  (
    .i0(\t/a/MEM_aludat [19]),
    .i1(\t/a/memreaddat [19]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [19]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b2  (
    .i0(\t/a/MEM_aludat [2]),
    .i1(\t/a/memreaddat [2]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [2]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b20  (
    .i0(\t/a/MEM_aludat [20]),
    .i1(\t/a/memreaddat [20]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [20]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b21  (
    .i0(\t/a/MEM_aludat [21]),
    .i1(\t/a/memreaddat [21]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [21]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b22  (
    .i0(\t/a/MEM_aludat [22]),
    .i1(\t/a/memreaddat [22]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [22]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b23  (
    .i0(\t/a/MEM_aludat [23]),
    .i1(\t/a/memreaddat [23]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [23]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b24  (
    .i0(\t/a/MEM_aludat [24]),
    .i1(\t/a/memreaddat [24]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [24]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b25  (
    .i0(\t/a/MEM_aludat [25]),
    .i1(\t/a/memreaddat [25]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [25]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b26  (
    .i0(\t/a/MEM_aludat [26]),
    .i1(\t/a/memreaddat [26]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [26]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b27  (
    .i0(\t/a/MEM_aludat [27]),
    .i1(\t/a/memreaddat [27]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [27]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b28  (
    .i0(\t/a/MEM_aludat [28]),
    .i1(\t/a/memreaddat [28]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [28]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b29  (
    .i0(\t/a/MEM_aludat [29]),
    .i1(\t/a/memreaddat [29]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [29]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b3  (
    .i0(\t/a/MEM_aludat [3]),
    .i1(\t/a/memreaddat [3]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [3]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b30  (
    .i0(\t/a/MEM_aludat [30]),
    .i1(\t/a/memreaddat [30]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [30]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b31  (
    .i0(\t/a/MEM_aludat [31]),
    .i1(\t/a/memreaddat [31]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [31]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b4  (
    .i0(\t/a/MEM_aludat [4]),
    .i1(\t/a/memreaddat [4]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [4]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b5  (
    .i0(\t/a/MEM_aludat [5]),
    .i1(\t/a/memreaddat [5]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [5]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b6  (
    .i0(\t/a/MEM_aludat [6]),
    .i1(\t/a/memreaddat [6]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [6]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b7  (
    .i0(\t/a/MEM_aludat [7]),
    .i1(\t/a/memreaddat [7]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [7]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b8  (
    .i0(\t/a/MEM_aludat [8]),
    .i1(\t/a/memreaddat [8]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [8]));  // flow_line_reg.v(227)
  binary_mux_s1_w1 \t/a/mem_wb/mux0_b9  (
    .i0(\t/a/MEM_aludat [9]),
    .i1(\t/a/memreaddat [9]),
    .sel(\t/memread_cs ),
    .o(\t/a/mem_wb/n5 [9]));  // flow_line_reg.v(227)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b0  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [0]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b1  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [1]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b10  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [10]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [10]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b11  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [11]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [11]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b12  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [12]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [12]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b13  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [13]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [13]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b14  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [14]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [14]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b15  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [15]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [15]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b16  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [16]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [16]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b17  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [17]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [17]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b18  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [18]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [18]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b19  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [19]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [19]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b2  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [2]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b20  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [20]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [20]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b21  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [21]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [21]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b22  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [22]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [22]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b23  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [23]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [23]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b24  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [24]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [24]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b25  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [25]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [25]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b26  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [26]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [26]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b27  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [27]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [27]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b28  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [28]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [28]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b29  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [29]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [29]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b3  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [3]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b30  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [30]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [30]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b31  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [31]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [31]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b4  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [4]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b5  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [5]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [5]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b6  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [6]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [6]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b7  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [7]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [7]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b8  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [8]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [8]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg0_b9  (
    .clk(clock),
    .d(\t/a/mem_wb/n5 [9]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/reg_writedat [9]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg1_b0  (
    .clk(clock),
    .d(\t/a/MEM_op [0]),
    .en(~\t/a/ex_mem/n0 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\t/a/WB_op [0]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg1_b1  (
    .clk(clock),
    .d(\t/a/MEM_op [1]),
    .en(~\t/a/ex_mem/n0 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\t/a/WB_op [1]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg1_b2  (
    .clk(clock),
    .d(\t/a/MEM_op [2]),
    .en(~\t/a/ex_mem/n0 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\t/a/WB_op [2]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg1_b3  (
    .clk(clock),
    .d(\t/a/MEM_op [3]),
    .en(~\t/a/ex_mem/n0 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\t/a/WB_op [3]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg1_b4  (
    .clk(clock),
    .d(\t/a/MEM_op [4]),
    .en(~\t/a/ex_mem/n0 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\t/a/WB_op [4]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg1_b5  (
    .clk(clock),
    .d(\t/a/MEM_op [5]),
    .en(~\t/a/ex_mem/n0 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\t/a/WB_op [5]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg1_b6  (
    .clk(clock),
    .d(\t/a/MEM_op [6]),
    .en(~\t/a/ex_mem/n0 ),
    .reset(1'b0),
    .set(1'b0),
    .q(\t/a/WB_op [6]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg2_b0  (
    .clk(clock),
    .d(\t/a/MEM_rd [0]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/WB_rd [0]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg2_b1  (
    .clk(clock),
    .d(\t/a/MEM_rd [1]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/WB_rd [1]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg2_b2  (
    .clk(clock),
    .d(\t/a/MEM_rd [2]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/WB_rd [2]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg2_b3  (
    .clk(clock),
    .d(\t/a/MEM_rd [3]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/WB_rd [3]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/reg2_b4  (
    .clk(clock),
    .d(\t/a/MEM_rd [4]),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/WB_rd [4]));  // flow_line_reg.v(234)
  reg_ar_as_w1 \t/a/mem_wb/regwritecs_reg  (
    .clk(clock),
    .d(\t/a/mem_wb/n12 ),
    .en(1'b1),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/WB_regwritecs ));  // flow_line_reg.v(234)
  or \t/a/mem_wb/u10  (\t/a/mem_wb/n10 , \t/a/mem_wb/n8 , \t/a/mem_wb/n9 );  // flow_line_reg.v(230)
  AL_MUX \t/a/mem_wb/u12  (
    .i0(\t/a/mem_wb/n11 ),
    .i1(1'b0),
    .sel(\t/a/mem_wb/n10 ),
    .o(\t/a/mem_wb/n12 ));  // flow_line_reg.v(233)
  or \t/a/mem_wb/u13  (\t/a/mem_wb/n14 , \t/a/MEM_op [5], \t/a/MEM_op [6]);  // flow_line_reg.v(232)
  or \t/a/mem_wb/u14  (\t/a/mem_wb/n13 , \t/a/mem_wb/n0 , \t/a/mem_wb/n14 );  // flow_line_reg.v(232)
  or \t/a/mem_wb/u15  (\t/a/mem_wb/n11 , \t/a/mem_wb/n1 , \t/a/mem_wb/n13 );  // flow_line_reg.v(232)
  or \t/a/mem_wb/u2  (\t/a/mem_wb/n0 , \t/a/MEM_op [3], \t/a/MEM_op [4]);  // flow_line_reg.v(232)
  or \t/a/mem_wb/u3  (\t/a/mem_wb/n1 , \t/a/MEM_op [0], \t/a/mem_wb/n2 );  // flow_line_reg.v(232)
  or \t/a/mem_wb/u7  (\t/a/mem_wb/n2 , \t/a/MEM_op [1], \t/a/MEM_op [2]);  // flow_line_reg.v(232)
  or \t/a/mem_wb/u9  (\t/a/mem_wb/n8 , memwrite_cs, \t/a/mem_wb/n7 );  // flow_line_reg.v(229)
  binary_mux_s1_w1 \t/a/mux0_b0  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\t/a/n14 ),
    .o(\t/a/alu_A_select [0]));  // cpu.v(249)
  binary_mux_s1_w1 \t/a/mux0_b1  (
    .i0(\t/a/n23 ),
    .i1(1'b0),
    .sel(\t/a/n14 ),
    .o(\t/a/alu_A_select [1]));  // cpu.v(249)
  binary_mux_s1_w1 \t/a/mux1_b0  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\t/a/n27 ),
    .o(\t/a/alu_B_select [0]));  // cpu.v(266)
  binary_mux_s1_w1 \t/a/mux1_b1  (
    .i0(\t/a/n31 ),
    .i1(1'b0),
    .sel(\t/a/n27 ),
    .o(\t/a/alu_B_select [1]));  // cpu.v(266)
  binary_mux_s1_w1 \t/a/mux2_b0  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [0]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [0]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b1  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [1]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [1]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b10  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [10]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [10]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b11  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [11]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [11]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b12  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [12]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [12]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b13  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [13]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [13]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b14  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [14]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [14]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b15  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [15]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [15]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b16  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [16]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [16]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b17  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [17]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [17]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b18  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [18]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [18]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b19  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [19]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [19]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b2  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [2]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [2]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b20  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [20]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [20]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b21  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [21]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [21]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b22  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [22]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [22]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b23  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [23]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [23]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b24  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [24]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [24]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b25  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [25]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [25]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b26  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [26]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [26]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b27  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [27]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [27]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b28  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [28]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [28]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b29  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [29]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [29]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b3  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [3]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [3]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b30  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [30]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [30]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b31  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [31]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [31]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b4  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [4]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [4]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b5  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [5]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [5]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b6  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [6]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [6]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b7  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [7]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [7]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b8  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [8]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [8]));  // cpu.v(290)
  binary_mux_s1_w1 \t/a/mux2_b9  (
    .i0(1'b0),
    .i1(\t/a/MEM_aludat [9]),
    .sel(\t/a/n34 ),
    .o(\t/memaddress [9]));  // cpu.v(290)
  and \t/a/mux3_b0_sel_is_1  (\t/a/mux3_b0_sel_is_1_o , memwrite_cs, \t/a/n33 );
  and \t/a/mux3_b10_sel_is_3  (\t/a/mux3_b10_sel_is_3_o , memwrite_cs, \t/a/sel0_b10_sel_o );
  and \t/a/mux3_b16_sel_is_3  (\t/a/mux3_b16_sel_is_3_o , memwrite_cs, \t/a/n37 );
  binary_mux_s3_w1 \t/a/mux4_b0  (
    .i0(\t/memreaddat [0]),
    .i1(\t/memreaddat [0]),
    .i2(\t/memreaddat [0]),
    .i3(1'b0),
    .i4(\t/memreaddat [0]),
    .i5(\t/memreaddat [0]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [0]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b1  (
    .i0(\t/memreaddat [1]),
    .i1(\t/memreaddat [1]),
    .i2(\t/memreaddat [1]),
    .i3(1'b0),
    .i4(\t/memreaddat [1]),
    .i5(\t/memreaddat [1]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [1]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b10  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [10]),
    .i2(\t/memreaddat [10]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(\t/memreaddat [10]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [10]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b11  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [11]),
    .i2(\t/memreaddat [11]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(\t/memreaddat [11]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [11]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b12  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [12]),
    .i2(\t/memreaddat [12]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(\t/memreaddat [12]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [12]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b13  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [13]),
    .i2(\t/memreaddat [13]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(\t/memreaddat [13]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [13]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b14  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [14]),
    .i2(\t/memreaddat [14]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(\t/memreaddat [14]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [14]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b15  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [15]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(\t/memreaddat [15]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [15]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b16  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [16]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [16]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b17  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [17]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [17]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b18  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [18]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [18]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b19  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [19]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [19]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b2  (
    .i0(\t/memreaddat [2]),
    .i1(\t/memreaddat [2]),
    .i2(\t/memreaddat [2]),
    .i3(1'b0),
    .i4(\t/memreaddat [2]),
    .i5(\t/memreaddat [2]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [2]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b20  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [20]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [20]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b21  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [21]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [21]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b22  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [22]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [22]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b23  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [23]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [23]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b24  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [24]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [24]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b25  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [25]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [25]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b26  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [26]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [26]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b27  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [27]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [27]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b28  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [28]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [28]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b29  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [29]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [29]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b3  (
    .i0(\t/memreaddat [3]),
    .i1(\t/memreaddat [3]),
    .i2(\t/memreaddat [3]),
    .i3(1'b0),
    .i4(\t/memreaddat [3]),
    .i5(\t/memreaddat [3]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [3]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b30  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [30]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [30]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b31  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [15]),
    .i2(\t/memreaddat [31]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(1'b0),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [31]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b4  (
    .i0(\t/memreaddat [4]),
    .i1(\t/memreaddat [4]),
    .i2(\t/memreaddat [4]),
    .i3(1'b0),
    .i4(\t/memreaddat [4]),
    .i5(\t/memreaddat [4]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [4]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b5  (
    .i0(\t/memreaddat [5]),
    .i1(\t/memreaddat [5]),
    .i2(\t/memreaddat [5]),
    .i3(1'b0),
    .i4(\t/memreaddat [5]),
    .i5(\t/memreaddat [5]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [5]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b6  (
    .i0(\t/memreaddat [6]),
    .i1(\t/memreaddat [6]),
    .i2(\t/memreaddat [6]),
    .i3(1'b0),
    .i4(\t/memreaddat [6]),
    .i5(\t/memreaddat [6]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [6]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b7  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [7]),
    .i2(\t/memreaddat [7]),
    .i3(1'b0),
    .i4(\t/memreaddat [7]),
    .i5(\t/memreaddat [7]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [7]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b8  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [8]),
    .i2(\t/memreaddat [8]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(\t/memreaddat [8]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [8]));  // cpu.v(320)
  binary_mux_s3_w1 \t/a/mux4_b9  (
    .i0(\t/memreaddat [7]),
    .i1(\t/memreaddat [9]),
    .i2(\t/memreaddat [9]),
    .i3(1'b0),
    .i4(1'b0),
    .i5(\t/memreaddat [9]),
    .i6(1'b0),
    .i7(1'b0),
    .sel(\t/a/MEM_fun3 ),
    .o(\t/a/n40 [9]));  // cpu.v(320)
  binary_mux_s1_w1 \t/a/mux5_b0  (
    .i0(1'b0),
    .i1(\t/a/n40 [0]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [0]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b1  (
    .i0(1'b0),
    .i1(\t/a/n40 [1]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [1]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b10  (
    .i0(1'b0),
    .i1(\t/a/n40 [10]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [10]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b11  (
    .i0(1'b0),
    .i1(\t/a/n40 [11]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [11]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b12  (
    .i0(1'b0),
    .i1(\t/a/n40 [12]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [12]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b13  (
    .i0(1'b0),
    .i1(\t/a/n40 [13]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [13]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b14  (
    .i0(1'b0),
    .i1(\t/a/n40 [14]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [14]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b15  (
    .i0(1'b0),
    .i1(\t/a/n40 [15]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [15]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b16  (
    .i0(1'b0),
    .i1(\t/a/n40 [16]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [16]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b17  (
    .i0(1'b0),
    .i1(\t/a/n40 [17]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [17]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b18  (
    .i0(1'b0),
    .i1(\t/a/n40 [18]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [18]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b19  (
    .i0(1'b0),
    .i1(\t/a/n40 [19]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [19]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b2  (
    .i0(1'b0),
    .i1(\t/a/n40 [2]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [2]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b20  (
    .i0(1'b0),
    .i1(\t/a/n40 [20]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [20]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b21  (
    .i0(1'b0),
    .i1(\t/a/n40 [21]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [21]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b22  (
    .i0(1'b0),
    .i1(\t/a/n40 [22]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [22]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b23  (
    .i0(1'b0),
    .i1(\t/a/n40 [23]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [23]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b24  (
    .i0(1'b0),
    .i1(\t/a/n40 [24]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [24]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b25  (
    .i0(1'b0),
    .i1(\t/a/n40 [25]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [25]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b26  (
    .i0(1'b0),
    .i1(\t/a/n40 [26]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [26]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b27  (
    .i0(1'b0),
    .i1(\t/a/n40 [27]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [27]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b28  (
    .i0(1'b0),
    .i1(\t/a/n40 [28]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [28]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b29  (
    .i0(1'b0),
    .i1(\t/a/n40 [29]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [29]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b3  (
    .i0(1'b0),
    .i1(\t/a/n40 [3]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [3]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b30  (
    .i0(1'b0),
    .i1(\t/a/n40 [30]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [30]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b31  (
    .i0(1'b0),
    .i1(\t/a/n40 [31]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [31]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b4  (
    .i0(1'b0),
    .i1(\t/a/n40 [4]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [4]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b5  (
    .i0(1'b0),
    .i1(\t/a/n40 [5]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [5]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b6  (
    .i0(1'b0),
    .i1(\t/a/n40 [6]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [6]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b7  (
    .i0(1'b0),
    .i1(\t/a/n40 [7]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [7]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b8  (
    .i0(1'b0),
    .i1(\t/a/n40 [8]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [8]));  // cpu.v(326)
  binary_mux_s1_w1 \t/a/mux5_b9  (
    .i0(1'b0),
    .i1(\t/a/n40 [9]),
    .sel(\t/memread_cs ),
    .o(\t/a/memreaddat [9]));  // cpu.v(326)
  ne_w7 \t/a/neq0  (
    .i0(\t/instruction [6:0]),
    .i1(7'b1100011),
    .o(\t/a/n1 ));  // cpu.v(179)
  ne_w7 \t/a/neq1  (
    .i0(\t/a/MEM_op ),
    .i1(7'b0100011),
    .o(\t/a/n6 ));  // cpu.v(237)
  ne_w7 \t/a/neq2  (
    .i0(\t/a/MEM_op ),
    .i1(7'b1100011),
    .o(\t/a/n7 ));  // cpu.v(238)
  ne_w5 \t/a/neq3  (
    .i0(\t/a/MEM_rd ),
    .i1(5'b00000),
    .o(\t/a/n11 ));  // cpu.v(240)
  ne_w7 \t/a/neq4  (
    .i0(\t/a/MEM_op ),
    .i1(7'b0000011),
    .o(\t/a/n13 ));  // cpu.v(241)
  ne_w7 \t/a/neq5  (
    .i0(\t/a/WB_op ),
    .i1(7'b0100011),
    .o(\t/a/n15 ));  // cpu.v(243)
  ne_w7 \t/a/neq6  (
    .i0(\t/a/WB_op ),
    .i1(7'b1100011),
    .o(\t/a/n16 ));  // cpu.v(244)
  ne_w5 \t/a/neq7  (
    .i0(\t/a/WB_rd ),
    .i1(5'b00000),
    .o(\t/a/n18 ));  // cpu.v(245)
  ne_w5 \t/a/neq8  (
    .i0(\t/a/MEM_rd ),
    .i1(\t/a/EX_rs1 ),
    .o(\t/a/n22 ));  // cpu.v(247)
  ne_w5 \t/a/neq9  (
    .i0(\t/a/MEM_rd ),
    .i1(\t/a/EX_rs2 ),
    .o(\t/a/n30 ));  // cpu.v(264)
  eq_w1 \t/a/regfile/eq0  (
    .i0(\t/a/WB_regwritecs ),
    .i1(1'b1),
    .o(\t/a/regfile/n0 ));  // register.v(10)
  eq_w5 \t/a/regfile/eq1  (
    .i0(\t/a/WB_rd ),
    .i1(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n1 ));  // register.v(10)
  eq_w5 \t/a/regfile/eq2  (
    .i0(\t/a/WB_rd ),
    .i1(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n3 ));  // register.v(10)
  binary_mux_s5_w1 \t/a/regfile/mux0_b0  (
    .i0(\t/a/regfile/regfile$0$ [0]),
    .i1(\t/a/regfile/regfile$1$ [0]),
    .i10(\t/a/regfile/regfile$10$ [0]),
    .i11(\t/a/regfile/regfile$11$ [0]),
    .i12(\t/a/regfile/regfile$12$ [0]),
    .i13(\t/a/regfile/regfile$13$ [0]),
    .i14(\t/a/regfile/regfile$14$ [0]),
    .i15(\t/a/regfile/regfile$15$ [0]),
    .i16(\t/a/regfile/regfile$16$ [0]),
    .i17(\t/a/regfile/regfile$17$ [0]),
    .i18(\t/a/regfile/regfile$18$ [0]),
    .i19(\t/a/regfile/regfile$19$ [0]),
    .i2(\t/a/regfile/regfile$2$ [0]),
    .i20(\t/a/regfile/regfile$20$ [0]),
    .i21(\t/a/regfile/regfile$21$ [0]),
    .i22(\t/a/regfile/regfile$22$ [0]),
    .i23(\t/a/regfile/regfile$23$ [0]),
    .i24(\t/a/regfile/regfile$24$ [0]),
    .i25(\t/a/regfile/regfile$25$ [0]),
    .i26(\t/a/regfile/regfile$26$ [0]),
    .i27(\t/a/regfile/regfile$27$ [0]),
    .i28(\t/a/regfile/regfile$28$ [0]),
    .i29(\t/a/regfile/regfile$29$ [0]),
    .i3(\t/a/regfile/regfile$3$ [0]),
    .i30(\t/a/regfile/regfile$30$ [0]),
    .i31(\t/a/regfile/regfile$31$ [0]),
    .i4(\t/a/regfile/regfile$4$ [0]),
    .i5(\t/a/regfile/regfile$5$ [0]),
    .i6(\t/a/regfile/regfile$6$ [0]),
    .i7(\t/a/regfile/regfile$7$ [0]),
    .i8(\t/a/regfile/regfile$8$ [0]),
    .i9(\t/a/regfile/regfile$9$ [0]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [0]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b1  (
    .i0(\t/a/regfile/regfile$0$ [1]),
    .i1(\t/a/regfile/regfile$1$ [1]),
    .i10(\t/a/regfile/regfile$10$ [1]),
    .i11(\t/a/regfile/regfile$11$ [1]),
    .i12(\t/a/regfile/regfile$12$ [1]),
    .i13(\t/a/regfile/regfile$13$ [1]),
    .i14(\t/a/regfile/regfile$14$ [1]),
    .i15(\t/a/regfile/regfile$15$ [1]),
    .i16(\t/a/regfile/regfile$16$ [1]),
    .i17(\t/a/regfile/regfile$17$ [1]),
    .i18(\t/a/regfile/regfile$18$ [1]),
    .i19(\t/a/regfile/regfile$19$ [1]),
    .i2(\t/a/regfile/regfile$2$ [1]),
    .i20(\t/a/regfile/regfile$20$ [1]),
    .i21(\t/a/regfile/regfile$21$ [1]),
    .i22(\t/a/regfile/regfile$22$ [1]),
    .i23(\t/a/regfile/regfile$23$ [1]),
    .i24(\t/a/regfile/regfile$24$ [1]),
    .i25(\t/a/regfile/regfile$25$ [1]),
    .i26(\t/a/regfile/regfile$26$ [1]),
    .i27(\t/a/regfile/regfile$27$ [1]),
    .i28(\t/a/regfile/regfile$28$ [1]),
    .i29(\t/a/regfile/regfile$29$ [1]),
    .i3(\t/a/regfile/regfile$3$ [1]),
    .i30(\t/a/regfile/regfile$30$ [1]),
    .i31(\t/a/regfile/regfile$31$ [1]),
    .i4(\t/a/regfile/regfile$4$ [1]),
    .i5(\t/a/regfile/regfile$5$ [1]),
    .i6(\t/a/regfile/regfile$6$ [1]),
    .i7(\t/a/regfile/regfile$7$ [1]),
    .i8(\t/a/regfile/regfile$8$ [1]),
    .i9(\t/a/regfile/regfile$9$ [1]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [1]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b10  (
    .i0(\t/a/regfile/regfile$0$ [10]),
    .i1(\t/a/regfile/regfile$1$ [10]),
    .i10(\t/a/regfile/regfile$10$ [10]),
    .i11(\t/a/regfile/regfile$11$ [10]),
    .i12(\t/a/regfile/regfile$12$ [10]),
    .i13(\t/a/regfile/regfile$13$ [10]),
    .i14(\t/a/regfile/regfile$14$ [10]),
    .i15(\t/a/regfile/regfile$15$ [10]),
    .i16(\t/a/regfile/regfile$16$ [10]),
    .i17(\t/a/regfile/regfile$17$ [10]),
    .i18(\t/a/regfile/regfile$18$ [10]),
    .i19(\t/a/regfile/regfile$19$ [10]),
    .i2(\t/a/regfile/regfile$2$ [10]),
    .i20(\t/a/regfile/regfile$20$ [10]),
    .i21(\t/a/regfile/regfile$21$ [10]),
    .i22(\t/a/regfile/regfile$22$ [10]),
    .i23(\t/a/regfile/regfile$23$ [10]),
    .i24(\t/a/regfile/regfile$24$ [10]),
    .i25(\t/a/regfile/regfile$25$ [10]),
    .i26(\t/a/regfile/regfile$26$ [10]),
    .i27(\t/a/regfile/regfile$27$ [10]),
    .i28(\t/a/regfile/regfile$28$ [10]),
    .i29(\t/a/regfile/regfile$29$ [10]),
    .i3(\t/a/regfile/regfile$3$ [10]),
    .i30(\t/a/regfile/regfile$30$ [10]),
    .i31(\t/a/regfile/regfile$31$ [10]),
    .i4(\t/a/regfile/regfile$4$ [10]),
    .i5(\t/a/regfile/regfile$5$ [10]),
    .i6(\t/a/regfile/regfile$6$ [10]),
    .i7(\t/a/regfile/regfile$7$ [10]),
    .i8(\t/a/regfile/regfile$8$ [10]),
    .i9(\t/a/regfile/regfile$9$ [10]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [10]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b11  (
    .i0(\t/a/regfile/regfile$0$ [11]),
    .i1(\t/a/regfile/regfile$1$ [11]),
    .i10(\t/a/regfile/regfile$10$ [11]),
    .i11(\t/a/regfile/regfile$11$ [11]),
    .i12(\t/a/regfile/regfile$12$ [11]),
    .i13(\t/a/regfile/regfile$13$ [11]),
    .i14(\t/a/regfile/regfile$14$ [11]),
    .i15(\t/a/regfile/regfile$15$ [11]),
    .i16(\t/a/regfile/regfile$16$ [11]),
    .i17(\t/a/regfile/regfile$17$ [11]),
    .i18(\t/a/regfile/regfile$18$ [11]),
    .i19(\t/a/regfile/regfile$19$ [11]),
    .i2(\t/a/regfile/regfile$2$ [11]),
    .i20(\t/a/regfile/regfile$20$ [11]),
    .i21(\t/a/regfile/regfile$21$ [11]),
    .i22(\t/a/regfile/regfile$22$ [11]),
    .i23(\t/a/regfile/regfile$23$ [11]),
    .i24(\t/a/regfile/regfile$24$ [11]),
    .i25(\t/a/regfile/regfile$25$ [11]),
    .i26(\t/a/regfile/regfile$26$ [11]),
    .i27(\t/a/regfile/regfile$27$ [11]),
    .i28(\t/a/regfile/regfile$28$ [11]),
    .i29(\t/a/regfile/regfile$29$ [11]),
    .i3(\t/a/regfile/regfile$3$ [11]),
    .i30(\t/a/regfile/regfile$30$ [11]),
    .i31(\t/a/regfile/regfile$31$ [11]),
    .i4(\t/a/regfile/regfile$4$ [11]),
    .i5(\t/a/regfile/regfile$5$ [11]),
    .i6(\t/a/regfile/regfile$6$ [11]),
    .i7(\t/a/regfile/regfile$7$ [11]),
    .i8(\t/a/regfile/regfile$8$ [11]),
    .i9(\t/a/regfile/regfile$9$ [11]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [11]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b12  (
    .i0(\t/a/regfile/regfile$0$ [12]),
    .i1(\t/a/regfile/regfile$1$ [12]),
    .i10(\t/a/regfile/regfile$10$ [12]),
    .i11(\t/a/regfile/regfile$11$ [12]),
    .i12(\t/a/regfile/regfile$12$ [12]),
    .i13(\t/a/regfile/regfile$13$ [12]),
    .i14(\t/a/regfile/regfile$14$ [12]),
    .i15(\t/a/regfile/regfile$15$ [12]),
    .i16(\t/a/regfile/regfile$16$ [12]),
    .i17(\t/a/regfile/regfile$17$ [12]),
    .i18(\t/a/regfile/regfile$18$ [12]),
    .i19(\t/a/regfile/regfile$19$ [12]),
    .i2(\t/a/regfile/regfile$2$ [12]),
    .i20(\t/a/regfile/regfile$20$ [12]),
    .i21(\t/a/regfile/regfile$21$ [12]),
    .i22(\t/a/regfile/regfile$22$ [12]),
    .i23(\t/a/regfile/regfile$23$ [12]),
    .i24(\t/a/regfile/regfile$24$ [12]),
    .i25(\t/a/regfile/regfile$25$ [12]),
    .i26(\t/a/regfile/regfile$26$ [12]),
    .i27(\t/a/regfile/regfile$27$ [12]),
    .i28(\t/a/regfile/regfile$28$ [12]),
    .i29(\t/a/regfile/regfile$29$ [12]),
    .i3(\t/a/regfile/regfile$3$ [12]),
    .i30(\t/a/regfile/regfile$30$ [12]),
    .i31(\t/a/regfile/regfile$31$ [12]),
    .i4(\t/a/regfile/regfile$4$ [12]),
    .i5(\t/a/regfile/regfile$5$ [12]),
    .i6(\t/a/regfile/regfile$6$ [12]),
    .i7(\t/a/regfile/regfile$7$ [12]),
    .i8(\t/a/regfile/regfile$8$ [12]),
    .i9(\t/a/regfile/regfile$9$ [12]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [12]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b13  (
    .i0(\t/a/regfile/regfile$0$ [13]),
    .i1(\t/a/regfile/regfile$1$ [13]),
    .i10(\t/a/regfile/regfile$10$ [13]),
    .i11(\t/a/regfile/regfile$11$ [13]),
    .i12(\t/a/regfile/regfile$12$ [13]),
    .i13(\t/a/regfile/regfile$13$ [13]),
    .i14(\t/a/regfile/regfile$14$ [13]),
    .i15(\t/a/regfile/regfile$15$ [13]),
    .i16(\t/a/regfile/regfile$16$ [13]),
    .i17(\t/a/regfile/regfile$17$ [13]),
    .i18(\t/a/regfile/regfile$18$ [13]),
    .i19(\t/a/regfile/regfile$19$ [13]),
    .i2(\t/a/regfile/regfile$2$ [13]),
    .i20(\t/a/regfile/regfile$20$ [13]),
    .i21(\t/a/regfile/regfile$21$ [13]),
    .i22(\t/a/regfile/regfile$22$ [13]),
    .i23(\t/a/regfile/regfile$23$ [13]),
    .i24(\t/a/regfile/regfile$24$ [13]),
    .i25(\t/a/regfile/regfile$25$ [13]),
    .i26(\t/a/regfile/regfile$26$ [13]),
    .i27(\t/a/regfile/regfile$27$ [13]),
    .i28(\t/a/regfile/regfile$28$ [13]),
    .i29(\t/a/regfile/regfile$29$ [13]),
    .i3(\t/a/regfile/regfile$3$ [13]),
    .i30(\t/a/regfile/regfile$30$ [13]),
    .i31(\t/a/regfile/regfile$31$ [13]),
    .i4(\t/a/regfile/regfile$4$ [13]),
    .i5(\t/a/regfile/regfile$5$ [13]),
    .i6(\t/a/regfile/regfile$6$ [13]),
    .i7(\t/a/regfile/regfile$7$ [13]),
    .i8(\t/a/regfile/regfile$8$ [13]),
    .i9(\t/a/regfile/regfile$9$ [13]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [13]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b14  (
    .i0(\t/a/regfile/regfile$0$ [14]),
    .i1(\t/a/regfile/regfile$1$ [14]),
    .i10(\t/a/regfile/regfile$10$ [14]),
    .i11(\t/a/regfile/regfile$11$ [14]),
    .i12(\t/a/regfile/regfile$12$ [14]),
    .i13(\t/a/regfile/regfile$13$ [14]),
    .i14(\t/a/regfile/regfile$14$ [14]),
    .i15(\t/a/regfile/regfile$15$ [14]),
    .i16(\t/a/regfile/regfile$16$ [14]),
    .i17(\t/a/regfile/regfile$17$ [14]),
    .i18(\t/a/regfile/regfile$18$ [14]),
    .i19(\t/a/regfile/regfile$19$ [14]),
    .i2(\t/a/regfile/regfile$2$ [14]),
    .i20(\t/a/regfile/regfile$20$ [14]),
    .i21(\t/a/regfile/regfile$21$ [14]),
    .i22(\t/a/regfile/regfile$22$ [14]),
    .i23(\t/a/regfile/regfile$23$ [14]),
    .i24(\t/a/regfile/regfile$24$ [14]),
    .i25(\t/a/regfile/regfile$25$ [14]),
    .i26(\t/a/regfile/regfile$26$ [14]),
    .i27(\t/a/regfile/regfile$27$ [14]),
    .i28(\t/a/regfile/regfile$28$ [14]),
    .i29(\t/a/regfile/regfile$29$ [14]),
    .i3(\t/a/regfile/regfile$3$ [14]),
    .i30(\t/a/regfile/regfile$30$ [14]),
    .i31(\t/a/regfile/regfile$31$ [14]),
    .i4(\t/a/regfile/regfile$4$ [14]),
    .i5(\t/a/regfile/regfile$5$ [14]),
    .i6(\t/a/regfile/regfile$6$ [14]),
    .i7(\t/a/regfile/regfile$7$ [14]),
    .i8(\t/a/regfile/regfile$8$ [14]),
    .i9(\t/a/regfile/regfile$9$ [14]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [14]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b15  (
    .i0(\t/a/regfile/regfile$0$ [15]),
    .i1(\t/a/regfile/regfile$1$ [15]),
    .i10(\t/a/regfile/regfile$10$ [15]),
    .i11(\t/a/regfile/regfile$11$ [15]),
    .i12(\t/a/regfile/regfile$12$ [15]),
    .i13(\t/a/regfile/regfile$13$ [15]),
    .i14(\t/a/regfile/regfile$14$ [15]),
    .i15(\t/a/regfile/regfile$15$ [15]),
    .i16(\t/a/regfile/regfile$16$ [15]),
    .i17(\t/a/regfile/regfile$17$ [15]),
    .i18(\t/a/regfile/regfile$18$ [15]),
    .i19(\t/a/regfile/regfile$19$ [15]),
    .i2(\t/a/regfile/regfile$2$ [15]),
    .i20(\t/a/regfile/regfile$20$ [15]),
    .i21(\t/a/regfile/regfile$21$ [15]),
    .i22(\t/a/regfile/regfile$22$ [15]),
    .i23(\t/a/regfile/regfile$23$ [15]),
    .i24(\t/a/regfile/regfile$24$ [15]),
    .i25(\t/a/regfile/regfile$25$ [15]),
    .i26(\t/a/regfile/regfile$26$ [15]),
    .i27(\t/a/regfile/regfile$27$ [15]),
    .i28(\t/a/regfile/regfile$28$ [15]),
    .i29(\t/a/regfile/regfile$29$ [15]),
    .i3(\t/a/regfile/regfile$3$ [15]),
    .i30(\t/a/regfile/regfile$30$ [15]),
    .i31(\t/a/regfile/regfile$31$ [15]),
    .i4(\t/a/regfile/regfile$4$ [15]),
    .i5(\t/a/regfile/regfile$5$ [15]),
    .i6(\t/a/regfile/regfile$6$ [15]),
    .i7(\t/a/regfile/regfile$7$ [15]),
    .i8(\t/a/regfile/regfile$8$ [15]),
    .i9(\t/a/regfile/regfile$9$ [15]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [15]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b16  (
    .i0(\t/a/regfile/regfile$0$ [16]),
    .i1(\t/a/regfile/regfile$1$ [16]),
    .i10(\t/a/regfile/regfile$10$ [16]),
    .i11(\t/a/regfile/regfile$11$ [16]),
    .i12(\t/a/regfile/regfile$12$ [16]),
    .i13(\t/a/regfile/regfile$13$ [16]),
    .i14(\t/a/regfile/regfile$14$ [16]),
    .i15(\t/a/regfile/regfile$15$ [16]),
    .i16(\t/a/regfile/regfile$16$ [16]),
    .i17(\t/a/regfile/regfile$17$ [16]),
    .i18(\t/a/regfile/regfile$18$ [16]),
    .i19(\t/a/regfile/regfile$19$ [16]),
    .i2(\t/a/regfile/regfile$2$ [16]),
    .i20(\t/a/regfile/regfile$20$ [16]),
    .i21(\t/a/regfile/regfile$21$ [16]),
    .i22(\t/a/regfile/regfile$22$ [16]),
    .i23(\t/a/regfile/regfile$23$ [16]),
    .i24(\t/a/regfile/regfile$24$ [16]),
    .i25(\t/a/regfile/regfile$25$ [16]),
    .i26(\t/a/regfile/regfile$26$ [16]),
    .i27(\t/a/regfile/regfile$27$ [16]),
    .i28(\t/a/regfile/regfile$28$ [16]),
    .i29(\t/a/regfile/regfile$29$ [16]),
    .i3(\t/a/regfile/regfile$3$ [16]),
    .i30(\t/a/regfile/regfile$30$ [16]),
    .i31(\t/a/regfile/regfile$31$ [16]),
    .i4(\t/a/regfile/regfile$4$ [16]),
    .i5(\t/a/regfile/regfile$5$ [16]),
    .i6(\t/a/regfile/regfile$6$ [16]),
    .i7(\t/a/regfile/regfile$7$ [16]),
    .i8(\t/a/regfile/regfile$8$ [16]),
    .i9(\t/a/regfile/regfile$9$ [16]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [16]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b17  (
    .i0(\t/a/regfile/regfile$0$ [17]),
    .i1(\t/a/regfile/regfile$1$ [17]),
    .i10(\t/a/regfile/regfile$10$ [17]),
    .i11(\t/a/regfile/regfile$11$ [17]),
    .i12(\t/a/regfile/regfile$12$ [17]),
    .i13(\t/a/regfile/regfile$13$ [17]),
    .i14(\t/a/regfile/regfile$14$ [17]),
    .i15(\t/a/regfile/regfile$15$ [17]),
    .i16(\t/a/regfile/regfile$16$ [17]),
    .i17(\t/a/regfile/regfile$17$ [17]),
    .i18(\t/a/regfile/regfile$18$ [17]),
    .i19(\t/a/regfile/regfile$19$ [17]),
    .i2(\t/a/regfile/regfile$2$ [17]),
    .i20(\t/a/regfile/regfile$20$ [17]),
    .i21(\t/a/regfile/regfile$21$ [17]),
    .i22(\t/a/regfile/regfile$22$ [17]),
    .i23(\t/a/regfile/regfile$23$ [17]),
    .i24(\t/a/regfile/regfile$24$ [17]),
    .i25(\t/a/regfile/regfile$25$ [17]),
    .i26(\t/a/regfile/regfile$26$ [17]),
    .i27(\t/a/regfile/regfile$27$ [17]),
    .i28(\t/a/regfile/regfile$28$ [17]),
    .i29(\t/a/regfile/regfile$29$ [17]),
    .i3(\t/a/regfile/regfile$3$ [17]),
    .i30(\t/a/regfile/regfile$30$ [17]),
    .i31(\t/a/regfile/regfile$31$ [17]),
    .i4(\t/a/regfile/regfile$4$ [17]),
    .i5(\t/a/regfile/regfile$5$ [17]),
    .i6(\t/a/regfile/regfile$6$ [17]),
    .i7(\t/a/regfile/regfile$7$ [17]),
    .i8(\t/a/regfile/regfile$8$ [17]),
    .i9(\t/a/regfile/regfile$9$ [17]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [17]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b18  (
    .i0(\t/a/regfile/regfile$0$ [18]),
    .i1(\t/a/regfile/regfile$1$ [18]),
    .i10(\t/a/regfile/regfile$10$ [18]),
    .i11(\t/a/regfile/regfile$11$ [18]),
    .i12(\t/a/regfile/regfile$12$ [18]),
    .i13(\t/a/regfile/regfile$13$ [18]),
    .i14(\t/a/regfile/regfile$14$ [18]),
    .i15(\t/a/regfile/regfile$15$ [18]),
    .i16(\t/a/regfile/regfile$16$ [18]),
    .i17(\t/a/regfile/regfile$17$ [18]),
    .i18(\t/a/regfile/regfile$18$ [18]),
    .i19(\t/a/regfile/regfile$19$ [18]),
    .i2(\t/a/regfile/regfile$2$ [18]),
    .i20(\t/a/regfile/regfile$20$ [18]),
    .i21(\t/a/regfile/regfile$21$ [18]),
    .i22(\t/a/regfile/regfile$22$ [18]),
    .i23(\t/a/regfile/regfile$23$ [18]),
    .i24(\t/a/regfile/regfile$24$ [18]),
    .i25(\t/a/regfile/regfile$25$ [18]),
    .i26(\t/a/regfile/regfile$26$ [18]),
    .i27(\t/a/regfile/regfile$27$ [18]),
    .i28(\t/a/regfile/regfile$28$ [18]),
    .i29(\t/a/regfile/regfile$29$ [18]),
    .i3(\t/a/regfile/regfile$3$ [18]),
    .i30(\t/a/regfile/regfile$30$ [18]),
    .i31(\t/a/regfile/regfile$31$ [18]),
    .i4(\t/a/regfile/regfile$4$ [18]),
    .i5(\t/a/regfile/regfile$5$ [18]),
    .i6(\t/a/regfile/regfile$6$ [18]),
    .i7(\t/a/regfile/regfile$7$ [18]),
    .i8(\t/a/regfile/regfile$8$ [18]),
    .i9(\t/a/regfile/regfile$9$ [18]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [18]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b19  (
    .i0(\t/a/regfile/regfile$0$ [19]),
    .i1(\t/a/regfile/regfile$1$ [19]),
    .i10(\t/a/regfile/regfile$10$ [19]),
    .i11(\t/a/regfile/regfile$11$ [19]),
    .i12(\t/a/regfile/regfile$12$ [19]),
    .i13(\t/a/regfile/regfile$13$ [19]),
    .i14(\t/a/regfile/regfile$14$ [19]),
    .i15(\t/a/regfile/regfile$15$ [19]),
    .i16(\t/a/regfile/regfile$16$ [19]),
    .i17(\t/a/regfile/regfile$17$ [19]),
    .i18(\t/a/regfile/regfile$18$ [19]),
    .i19(\t/a/regfile/regfile$19$ [19]),
    .i2(\t/a/regfile/regfile$2$ [19]),
    .i20(\t/a/regfile/regfile$20$ [19]),
    .i21(\t/a/regfile/regfile$21$ [19]),
    .i22(\t/a/regfile/regfile$22$ [19]),
    .i23(\t/a/regfile/regfile$23$ [19]),
    .i24(\t/a/regfile/regfile$24$ [19]),
    .i25(\t/a/regfile/regfile$25$ [19]),
    .i26(\t/a/regfile/regfile$26$ [19]),
    .i27(\t/a/regfile/regfile$27$ [19]),
    .i28(\t/a/regfile/regfile$28$ [19]),
    .i29(\t/a/regfile/regfile$29$ [19]),
    .i3(\t/a/regfile/regfile$3$ [19]),
    .i30(\t/a/regfile/regfile$30$ [19]),
    .i31(\t/a/regfile/regfile$31$ [19]),
    .i4(\t/a/regfile/regfile$4$ [19]),
    .i5(\t/a/regfile/regfile$5$ [19]),
    .i6(\t/a/regfile/regfile$6$ [19]),
    .i7(\t/a/regfile/regfile$7$ [19]),
    .i8(\t/a/regfile/regfile$8$ [19]),
    .i9(\t/a/regfile/regfile$9$ [19]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [19]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b2  (
    .i0(\t/a/regfile/regfile$0$ [2]),
    .i1(\t/a/regfile/regfile$1$ [2]),
    .i10(\t/a/regfile/regfile$10$ [2]),
    .i11(\t/a/regfile/regfile$11$ [2]),
    .i12(\t/a/regfile/regfile$12$ [2]),
    .i13(\t/a/regfile/regfile$13$ [2]),
    .i14(\t/a/regfile/regfile$14$ [2]),
    .i15(\t/a/regfile/regfile$15$ [2]),
    .i16(\t/a/regfile/regfile$16$ [2]),
    .i17(\t/a/regfile/regfile$17$ [2]),
    .i18(\t/a/regfile/regfile$18$ [2]),
    .i19(\t/a/regfile/regfile$19$ [2]),
    .i2(\t/a/regfile/regfile$2$ [2]),
    .i20(\t/a/regfile/regfile$20$ [2]),
    .i21(\t/a/regfile/regfile$21$ [2]),
    .i22(\t/a/regfile/regfile$22$ [2]),
    .i23(\t/a/regfile/regfile$23$ [2]),
    .i24(\t/a/regfile/regfile$24$ [2]),
    .i25(\t/a/regfile/regfile$25$ [2]),
    .i26(\t/a/regfile/regfile$26$ [2]),
    .i27(\t/a/regfile/regfile$27$ [2]),
    .i28(\t/a/regfile/regfile$28$ [2]),
    .i29(\t/a/regfile/regfile$29$ [2]),
    .i3(\t/a/regfile/regfile$3$ [2]),
    .i30(\t/a/regfile/regfile$30$ [2]),
    .i31(\t/a/regfile/regfile$31$ [2]),
    .i4(\t/a/regfile/regfile$4$ [2]),
    .i5(\t/a/regfile/regfile$5$ [2]),
    .i6(\t/a/regfile/regfile$6$ [2]),
    .i7(\t/a/regfile/regfile$7$ [2]),
    .i8(\t/a/regfile/regfile$8$ [2]),
    .i9(\t/a/regfile/regfile$9$ [2]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [2]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b20  (
    .i0(\t/a/regfile/regfile$0$ [20]),
    .i1(\t/a/regfile/regfile$1$ [20]),
    .i10(\t/a/regfile/regfile$10$ [20]),
    .i11(\t/a/regfile/regfile$11$ [20]),
    .i12(\t/a/regfile/regfile$12$ [20]),
    .i13(\t/a/regfile/regfile$13$ [20]),
    .i14(\t/a/regfile/regfile$14$ [20]),
    .i15(\t/a/regfile/regfile$15$ [20]),
    .i16(\t/a/regfile/regfile$16$ [20]),
    .i17(\t/a/regfile/regfile$17$ [20]),
    .i18(\t/a/regfile/regfile$18$ [20]),
    .i19(\t/a/regfile/regfile$19$ [20]),
    .i2(\t/a/regfile/regfile$2$ [20]),
    .i20(\t/a/regfile/regfile$20$ [20]),
    .i21(\t/a/regfile/regfile$21$ [20]),
    .i22(\t/a/regfile/regfile$22$ [20]),
    .i23(\t/a/regfile/regfile$23$ [20]),
    .i24(\t/a/regfile/regfile$24$ [20]),
    .i25(\t/a/regfile/regfile$25$ [20]),
    .i26(\t/a/regfile/regfile$26$ [20]),
    .i27(\t/a/regfile/regfile$27$ [20]),
    .i28(\t/a/regfile/regfile$28$ [20]),
    .i29(\t/a/regfile/regfile$29$ [20]),
    .i3(\t/a/regfile/regfile$3$ [20]),
    .i30(\t/a/regfile/regfile$30$ [20]),
    .i31(\t/a/regfile/regfile$31$ [20]),
    .i4(\t/a/regfile/regfile$4$ [20]),
    .i5(\t/a/regfile/regfile$5$ [20]),
    .i6(\t/a/regfile/regfile$6$ [20]),
    .i7(\t/a/regfile/regfile$7$ [20]),
    .i8(\t/a/regfile/regfile$8$ [20]),
    .i9(\t/a/regfile/regfile$9$ [20]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [20]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b21  (
    .i0(\t/a/regfile/regfile$0$ [21]),
    .i1(\t/a/regfile/regfile$1$ [21]),
    .i10(\t/a/regfile/regfile$10$ [21]),
    .i11(\t/a/regfile/regfile$11$ [21]),
    .i12(\t/a/regfile/regfile$12$ [21]),
    .i13(\t/a/regfile/regfile$13$ [21]),
    .i14(\t/a/regfile/regfile$14$ [21]),
    .i15(\t/a/regfile/regfile$15$ [21]),
    .i16(\t/a/regfile/regfile$16$ [21]),
    .i17(\t/a/regfile/regfile$17$ [21]),
    .i18(\t/a/regfile/regfile$18$ [21]),
    .i19(\t/a/regfile/regfile$19$ [21]),
    .i2(\t/a/regfile/regfile$2$ [21]),
    .i20(\t/a/regfile/regfile$20$ [21]),
    .i21(\t/a/regfile/regfile$21$ [21]),
    .i22(\t/a/regfile/regfile$22$ [21]),
    .i23(\t/a/regfile/regfile$23$ [21]),
    .i24(\t/a/regfile/regfile$24$ [21]),
    .i25(\t/a/regfile/regfile$25$ [21]),
    .i26(\t/a/regfile/regfile$26$ [21]),
    .i27(\t/a/regfile/regfile$27$ [21]),
    .i28(\t/a/regfile/regfile$28$ [21]),
    .i29(\t/a/regfile/regfile$29$ [21]),
    .i3(\t/a/regfile/regfile$3$ [21]),
    .i30(\t/a/regfile/regfile$30$ [21]),
    .i31(\t/a/regfile/regfile$31$ [21]),
    .i4(\t/a/regfile/regfile$4$ [21]),
    .i5(\t/a/regfile/regfile$5$ [21]),
    .i6(\t/a/regfile/regfile$6$ [21]),
    .i7(\t/a/regfile/regfile$7$ [21]),
    .i8(\t/a/regfile/regfile$8$ [21]),
    .i9(\t/a/regfile/regfile$9$ [21]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [21]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b22  (
    .i0(\t/a/regfile/regfile$0$ [22]),
    .i1(\t/a/regfile/regfile$1$ [22]),
    .i10(\t/a/regfile/regfile$10$ [22]),
    .i11(\t/a/regfile/regfile$11$ [22]),
    .i12(\t/a/regfile/regfile$12$ [22]),
    .i13(\t/a/regfile/regfile$13$ [22]),
    .i14(\t/a/regfile/regfile$14$ [22]),
    .i15(\t/a/regfile/regfile$15$ [22]),
    .i16(\t/a/regfile/regfile$16$ [22]),
    .i17(\t/a/regfile/regfile$17$ [22]),
    .i18(\t/a/regfile/regfile$18$ [22]),
    .i19(\t/a/regfile/regfile$19$ [22]),
    .i2(\t/a/regfile/regfile$2$ [22]),
    .i20(\t/a/regfile/regfile$20$ [22]),
    .i21(\t/a/regfile/regfile$21$ [22]),
    .i22(\t/a/regfile/regfile$22$ [22]),
    .i23(\t/a/regfile/regfile$23$ [22]),
    .i24(\t/a/regfile/regfile$24$ [22]),
    .i25(\t/a/regfile/regfile$25$ [22]),
    .i26(\t/a/regfile/regfile$26$ [22]),
    .i27(\t/a/regfile/regfile$27$ [22]),
    .i28(\t/a/regfile/regfile$28$ [22]),
    .i29(\t/a/regfile/regfile$29$ [22]),
    .i3(\t/a/regfile/regfile$3$ [22]),
    .i30(\t/a/regfile/regfile$30$ [22]),
    .i31(\t/a/regfile/regfile$31$ [22]),
    .i4(\t/a/regfile/regfile$4$ [22]),
    .i5(\t/a/regfile/regfile$5$ [22]),
    .i6(\t/a/regfile/regfile$6$ [22]),
    .i7(\t/a/regfile/regfile$7$ [22]),
    .i8(\t/a/regfile/regfile$8$ [22]),
    .i9(\t/a/regfile/regfile$9$ [22]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [22]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b23  (
    .i0(\t/a/regfile/regfile$0$ [23]),
    .i1(\t/a/regfile/regfile$1$ [23]),
    .i10(\t/a/regfile/regfile$10$ [23]),
    .i11(\t/a/regfile/regfile$11$ [23]),
    .i12(\t/a/regfile/regfile$12$ [23]),
    .i13(\t/a/regfile/regfile$13$ [23]),
    .i14(\t/a/regfile/regfile$14$ [23]),
    .i15(\t/a/regfile/regfile$15$ [23]),
    .i16(\t/a/regfile/regfile$16$ [23]),
    .i17(\t/a/regfile/regfile$17$ [23]),
    .i18(\t/a/regfile/regfile$18$ [23]),
    .i19(\t/a/regfile/regfile$19$ [23]),
    .i2(\t/a/regfile/regfile$2$ [23]),
    .i20(\t/a/regfile/regfile$20$ [23]),
    .i21(\t/a/regfile/regfile$21$ [23]),
    .i22(\t/a/regfile/regfile$22$ [23]),
    .i23(\t/a/regfile/regfile$23$ [23]),
    .i24(\t/a/regfile/regfile$24$ [23]),
    .i25(\t/a/regfile/regfile$25$ [23]),
    .i26(\t/a/regfile/regfile$26$ [23]),
    .i27(\t/a/regfile/regfile$27$ [23]),
    .i28(\t/a/regfile/regfile$28$ [23]),
    .i29(\t/a/regfile/regfile$29$ [23]),
    .i3(\t/a/regfile/regfile$3$ [23]),
    .i30(\t/a/regfile/regfile$30$ [23]),
    .i31(\t/a/regfile/regfile$31$ [23]),
    .i4(\t/a/regfile/regfile$4$ [23]),
    .i5(\t/a/regfile/regfile$5$ [23]),
    .i6(\t/a/regfile/regfile$6$ [23]),
    .i7(\t/a/regfile/regfile$7$ [23]),
    .i8(\t/a/regfile/regfile$8$ [23]),
    .i9(\t/a/regfile/regfile$9$ [23]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [23]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b24  (
    .i0(\t/a/regfile/regfile$0$ [24]),
    .i1(\t/a/regfile/regfile$1$ [24]),
    .i10(\t/a/regfile/regfile$10$ [24]),
    .i11(\t/a/regfile/regfile$11$ [24]),
    .i12(\t/a/regfile/regfile$12$ [24]),
    .i13(\t/a/regfile/regfile$13$ [24]),
    .i14(\t/a/regfile/regfile$14$ [24]),
    .i15(\t/a/regfile/regfile$15$ [24]),
    .i16(\t/a/regfile/regfile$16$ [24]),
    .i17(\t/a/regfile/regfile$17$ [24]),
    .i18(\t/a/regfile/regfile$18$ [24]),
    .i19(\t/a/regfile/regfile$19$ [24]),
    .i2(\t/a/regfile/regfile$2$ [24]),
    .i20(\t/a/regfile/regfile$20$ [24]),
    .i21(\t/a/regfile/regfile$21$ [24]),
    .i22(\t/a/regfile/regfile$22$ [24]),
    .i23(\t/a/regfile/regfile$23$ [24]),
    .i24(\t/a/regfile/regfile$24$ [24]),
    .i25(\t/a/regfile/regfile$25$ [24]),
    .i26(\t/a/regfile/regfile$26$ [24]),
    .i27(\t/a/regfile/regfile$27$ [24]),
    .i28(\t/a/regfile/regfile$28$ [24]),
    .i29(\t/a/regfile/regfile$29$ [24]),
    .i3(\t/a/regfile/regfile$3$ [24]),
    .i30(\t/a/regfile/regfile$30$ [24]),
    .i31(\t/a/regfile/regfile$31$ [24]),
    .i4(\t/a/regfile/regfile$4$ [24]),
    .i5(\t/a/regfile/regfile$5$ [24]),
    .i6(\t/a/regfile/regfile$6$ [24]),
    .i7(\t/a/regfile/regfile$7$ [24]),
    .i8(\t/a/regfile/regfile$8$ [24]),
    .i9(\t/a/regfile/regfile$9$ [24]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [24]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b25  (
    .i0(\t/a/regfile/regfile$0$ [25]),
    .i1(\t/a/regfile/regfile$1$ [25]),
    .i10(\t/a/regfile/regfile$10$ [25]),
    .i11(\t/a/regfile/regfile$11$ [25]),
    .i12(\t/a/regfile/regfile$12$ [25]),
    .i13(\t/a/regfile/regfile$13$ [25]),
    .i14(\t/a/regfile/regfile$14$ [25]),
    .i15(\t/a/regfile/regfile$15$ [25]),
    .i16(\t/a/regfile/regfile$16$ [25]),
    .i17(\t/a/regfile/regfile$17$ [25]),
    .i18(\t/a/regfile/regfile$18$ [25]),
    .i19(\t/a/regfile/regfile$19$ [25]),
    .i2(\t/a/regfile/regfile$2$ [25]),
    .i20(\t/a/regfile/regfile$20$ [25]),
    .i21(\t/a/regfile/regfile$21$ [25]),
    .i22(\t/a/regfile/regfile$22$ [25]),
    .i23(\t/a/regfile/regfile$23$ [25]),
    .i24(\t/a/regfile/regfile$24$ [25]),
    .i25(\t/a/regfile/regfile$25$ [25]),
    .i26(\t/a/regfile/regfile$26$ [25]),
    .i27(\t/a/regfile/regfile$27$ [25]),
    .i28(\t/a/regfile/regfile$28$ [25]),
    .i29(\t/a/regfile/regfile$29$ [25]),
    .i3(\t/a/regfile/regfile$3$ [25]),
    .i30(\t/a/regfile/regfile$30$ [25]),
    .i31(\t/a/regfile/regfile$31$ [25]),
    .i4(\t/a/regfile/regfile$4$ [25]),
    .i5(\t/a/regfile/regfile$5$ [25]),
    .i6(\t/a/regfile/regfile$6$ [25]),
    .i7(\t/a/regfile/regfile$7$ [25]),
    .i8(\t/a/regfile/regfile$8$ [25]),
    .i9(\t/a/regfile/regfile$9$ [25]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [25]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b26  (
    .i0(\t/a/regfile/regfile$0$ [26]),
    .i1(\t/a/regfile/regfile$1$ [26]),
    .i10(\t/a/regfile/regfile$10$ [26]),
    .i11(\t/a/regfile/regfile$11$ [26]),
    .i12(\t/a/regfile/regfile$12$ [26]),
    .i13(\t/a/regfile/regfile$13$ [26]),
    .i14(\t/a/regfile/regfile$14$ [26]),
    .i15(\t/a/regfile/regfile$15$ [26]),
    .i16(\t/a/regfile/regfile$16$ [26]),
    .i17(\t/a/regfile/regfile$17$ [26]),
    .i18(\t/a/regfile/regfile$18$ [26]),
    .i19(\t/a/regfile/regfile$19$ [26]),
    .i2(\t/a/regfile/regfile$2$ [26]),
    .i20(\t/a/regfile/regfile$20$ [26]),
    .i21(\t/a/regfile/regfile$21$ [26]),
    .i22(\t/a/regfile/regfile$22$ [26]),
    .i23(\t/a/regfile/regfile$23$ [26]),
    .i24(\t/a/regfile/regfile$24$ [26]),
    .i25(\t/a/regfile/regfile$25$ [26]),
    .i26(\t/a/regfile/regfile$26$ [26]),
    .i27(\t/a/regfile/regfile$27$ [26]),
    .i28(\t/a/regfile/regfile$28$ [26]),
    .i29(\t/a/regfile/regfile$29$ [26]),
    .i3(\t/a/regfile/regfile$3$ [26]),
    .i30(\t/a/regfile/regfile$30$ [26]),
    .i31(\t/a/regfile/regfile$31$ [26]),
    .i4(\t/a/regfile/regfile$4$ [26]),
    .i5(\t/a/regfile/regfile$5$ [26]),
    .i6(\t/a/regfile/regfile$6$ [26]),
    .i7(\t/a/regfile/regfile$7$ [26]),
    .i8(\t/a/regfile/regfile$8$ [26]),
    .i9(\t/a/regfile/regfile$9$ [26]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [26]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b27  (
    .i0(\t/a/regfile/regfile$0$ [27]),
    .i1(\t/a/regfile/regfile$1$ [27]),
    .i10(\t/a/regfile/regfile$10$ [27]),
    .i11(\t/a/regfile/regfile$11$ [27]),
    .i12(\t/a/regfile/regfile$12$ [27]),
    .i13(\t/a/regfile/regfile$13$ [27]),
    .i14(\t/a/regfile/regfile$14$ [27]),
    .i15(\t/a/regfile/regfile$15$ [27]),
    .i16(\t/a/regfile/regfile$16$ [27]),
    .i17(\t/a/regfile/regfile$17$ [27]),
    .i18(\t/a/regfile/regfile$18$ [27]),
    .i19(\t/a/regfile/regfile$19$ [27]),
    .i2(\t/a/regfile/regfile$2$ [27]),
    .i20(\t/a/regfile/regfile$20$ [27]),
    .i21(\t/a/regfile/regfile$21$ [27]),
    .i22(\t/a/regfile/regfile$22$ [27]),
    .i23(\t/a/regfile/regfile$23$ [27]),
    .i24(\t/a/regfile/regfile$24$ [27]),
    .i25(\t/a/regfile/regfile$25$ [27]),
    .i26(\t/a/regfile/regfile$26$ [27]),
    .i27(\t/a/regfile/regfile$27$ [27]),
    .i28(\t/a/regfile/regfile$28$ [27]),
    .i29(\t/a/regfile/regfile$29$ [27]),
    .i3(\t/a/regfile/regfile$3$ [27]),
    .i30(\t/a/regfile/regfile$30$ [27]),
    .i31(\t/a/regfile/regfile$31$ [27]),
    .i4(\t/a/regfile/regfile$4$ [27]),
    .i5(\t/a/regfile/regfile$5$ [27]),
    .i6(\t/a/regfile/regfile$6$ [27]),
    .i7(\t/a/regfile/regfile$7$ [27]),
    .i8(\t/a/regfile/regfile$8$ [27]),
    .i9(\t/a/regfile/regfile$9$ [27]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [27]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b28  (
    .i0(\t/a/regfile/regfile$0$ [28]),
    .i1(\t/a/regfile/regfile$1$ [28]),
    .i10(\t/a/regfile/regfile$10$ [28]),
    .i11(\t/a/regfile/regfile$11$ [28]),
    .i12(\t/a/regfile/regfile$12$ [28]),
    .i13(\t/a/regfile/regfile$13$ [28]),
    .i14(\t/a/regfile/regfile$14$ [28]),
    .i15(\t/a/regfile/regfile$15$ [28]),
    .i16(\t/a/regfile/regfile$16$ [28]),
    .i17(\t/a/regfile/regfile$17$ [28]),
    .i18(\t/a/regfile/regfile$18$ [28]),
    .i19(\t/a/regfile/regfile$19$ [28]),
    .i2(\t/a/regfile/regfile$2$ [28]),
    .i20(\t/a/regfile/regfile$20$ [28]),
    .i21(\t/a/regfile/regfile$21$ [28]),
    .i22(\t/a/regfile/regfile$22$ [28]),
    .i23(\t/a/regfile/regfile$23$ [28]),
    .i24(\t/a/regfile/regfile$24$ [28]),
    .i25(\t/a/regfile/regfile$25$ [28]),
    .i26(\t/a/regfile/regfile$26$ [28]),
    .i27(\t/a/regfile/regfile$27$ [28]),
    .i28(\t/a/regfile/regfile$28$ [28]),
    .i29(\t/a/regfile/regfile$29$ [28]),
    .i3(\t/a/regfile/regfile$3$ [28]),
    .i30(\t/a/regfile/regfile$30$ [28]),
    .i31(\t/a/regfile/regfile$31$ [28]),
    .i4(\t/a/regfile/regfile$4$ [28]),
    .i5(\t/a/regfile/regfile$5$ [28]),
    .i6(\t/a/regfile/regfile$6$ [28]),
    .i7(\t/a/regfile/regfile$7$ [28]),
    .i8(\t/a/regfile/regfile$8$ [28]),
    .i9(\t/a/regfile/regfile$9$ [28]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [28]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b29  (
    .i0(\t/a/regfile/regfile$0$ [29]),
    .i1(\t/a/regfile/regfile$1$ [29]),
    .i10(\t/a/regfile/regfile$10$ [29]),
    .i11(\t/a/regfile/regfile$11$ [29]),
    .i12(\t/a/regfile/regfile$12$ [29]),
    .i13(\t/a/regfile/regfile$13$ [29]),
    .i14(\t/a/regfile/regfile$14$ [29]),
    .i15(\t/a/regfile/regfile$15$ [29]),
    .i16(\t/a/regfile/regfile$16$ [29]),
    .i17(\t/a/regfile/regfile$17$ [29]),
    .i18(\t/a/regfile/regfile$18$ [29]),
    .i19(\t/a/regfile/regfile$19$ [29]),
    .i2(\t/a/regfile/regfile$2$ [29]),
    .i20(\t/a/regfile/regfile$20$ [29]),
    .i21(\t/a/regfile/regfile$21$ [29]),
    .i22(\t/a/regfile/regfile$22$ [29]),
    .i23(\t/a/regfile/regfile$23$ [29]),
    .i24(\t/a/regfile/regfile$24$ [29]),
    .i25(\t/a/regfile/regfile$25$ [29]),
    .i26(\t/a/regfile/regfile$26$ [29]),
    .i27(\t/a/regfile/regfile$27$ [29]),
    .i28(\t/a/regfile/regfile$28$ [29]),
    .i29(\t/a/regfile/regfile$29$ [29]),
    .i3(\t/a/regfile/regfile$3$ [29]),
    .i30(\t/a/regfile/regfile$30$ [29]),
    .i31(\t/a/regfile/regfile$31$ [29]),
    .i4(\t/a/regfile/regfile$4$ [29]),
    .i5(\t/a/regfile/regfile$5$ [29]),
    .i6(\t/a/regfile/regfile$6$ [29]),
    .i7(\t/a/regfile/regfile$7$ [29]),
    .i8(\t/a/regfile/regfile$8$ [29]),
    .i9(\t/a/regfile/regfile$9$ [29]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [29]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b3  (
    .i0(\t/a/regfile/regfile$0$ [3]),
    .i1(\t/a/regfile/regfile$1$ [3]),
    .i10(\t/a/regfile/regfile$10$ [3]),
    .i11(\t/a/regfile/regfile$11$ [3]),
    .i12(\t/a/regfile/regfile$12$ [3]),
    .i13(\t/a/regfile/regfile$13$ [3]),
    .i14(\t/a/regfile/regfile$14$ [3]),
    .i15(\t/a/regfile/regfile$15$ [3]),
    .i16(\t/a/regfile/regfile$16$ [3]),
    .i17(\t/a/regfile/regfile$17$ [3]),
    .i18(\t/a/regfile/regfile$18$ [3]),
    .i19(\t/a/regfile/regfile$19$ [3]),
    .i2(\t/a/regfile/regfile$2$ [3]),
    .i20(\t/a/regfile/regfile$20$ [3]),
    .i21(\t/a/regfile/regfile$21$ [3]),
    .i22(\t/a/regfile/regfile$22$ [3]),
    .i23(\t/a/regfile/regfile$23$ [3]),
    .i24(\t/a/regfile/regfile$24$ [3]),
    .i25(\t/a/regfile/regfile$25$ [3]),
    .i26(\t/a/regfile/regfile$26$ [3]),
    .i27(\t/a/regfile/regfile$27$ [3]),
    .i28(\t/a/regfile/regfile$28$ [3]),
    .i29(\t/a/regfile/regfile$29$ [3]),
    .i3(\t/a/regfile/regfile$3$ [3]),
    .i30(\t/a/regfile/regfile$30$ [3]),
    .i31(\t/a/regfile/regfile$31$ [3]),
    .i4(\t/a/regfile/regfile$4$ [3]),
    .i5(\t/a/regfile/regfile$5$ [3]),
    .i6(\t/a/regfile/regfile$6$ [3]),
    .i7(\t/a/regfile/regfile$7$ [3]),
    .i8(\t/a/regfile/regfile$8$ [3]),
    .i9(\t/a/regfile/regfile$9$ [3]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [3]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b30  (
    .i0(\t/a/regfile/regfile$0$ [30]),
    .i1(\t/a/regfile/regfile$1$ [30]),
    .i10(\t/a/regfile/regfile$10$ [30]),
    .i11(\t/a/regfile/regfile$11$ [30]),
    .i12(\t/a/regfile/regfile$12$ [30]),
    .i13(\t/a/regfile/regfile$13$ [30]),
    .i14(\t/a/regfile/regfile$14$ [30]),
    .i15(\t/a/regfile/regfile$15$ [30]),
    .i16(\t/a/regfile/regfile$16$ [30]),
    .i17(\t/a/regfile/regfile$17$ [30]),
    .i18(\t/a/regfile/regfile$18$ [30]),
    .i19(\t/a/regfile/regfile$19$ [30]),
    .i2(\t/a/regfile/regfile$2$ [30]),
    .i20(\t/a/regfile/regfile$20$ [30]),
    .i21(\t/a/regfile/regfile$21$ [30]),
    .i22(\t/a/regfile/regfile$22$ [30]),
    .i23(\t/a/regfile/regfile$23$ [30]),
    .i24(\t/a/regfile/regfile$24$ [30]),
    .i25(\t/a/regfile/regfile$25$ [30]),
    .i26(\t/a/regfile/regfile$26$ [30]),
    .i27(\t/a/regfile/regfile$27$ [30]),
    .i28(\t/a/regfile/regfile$28$ [30]),
    .i29(\t/a/regfile/regfile$29$ [30]),
    .i3(\t/a/regfile/regfile$3$ [30]),
    .i30(\t/a/regfile/regfile$30$ [30]),
    .i31(\t/a/regfile/regfile$31$ [30]),
    .i4(\t/a/regfile/regfile$4$ [30]),
    .i5(\t/a/regfile/regfile$5$ [30]),
    .i6(\t/a/regfile/regfile$6$ [30]),
    .i7(\t/a/regfile/regfile$7$ [30]),
    .i8(\t/a/regfile/regfile$8$ [30]),
    .i9(\t/a/regfile/regfile$9$ [30]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [30]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b31  (
    .i0(\t/a/regfile/regfile$0$ [31]),
    .i1(\t/a/regfile/regfile$1$ [31]),
    .i10(\t/a/regfile/regfile$10$ [31]),
    .i11(\t/a/regfile/regfile$11$ [31]),
    .i12(\t/a/regfile/regfile$12$ [31]),
    .i13(\t/a/regfile/regfile$13$ [31]),
    .i14(\t/a/regfile/regfile$14$ [31]),
    .i15(\t/a/regfile/regfile$15$ [31]),
    .i16(\t/a/regfile/regfile$16$ [31]),
    .i17(\t/a/regfile/regfile$17$ [31]),
    .i18(\t/a/regfile/regfile$18$ [31]),
    .i19(\t/a/regfile/regfile$19$ [31]),
    .i2(\t/a/regfile/regfile$2$ [31]),
    .i20(\t/a/regfile/regfile$20$ [31]),
    .i21(\t/a/regfile/regfile$21$ [31]),
    .i22(\t/a/regfile/regfile$22$ [31]),
    .i23(\t/a/regfile/regfile$23$ [31]),
    .i24(\t/a/regfile/regfile$24$ [31]),
    .i25(\t/a/regfile/regfile$25$ [31]),
    .i26(\t/a/regfile/regfile$26$ [31]),
    .i27(\t/a/regfile/regfile$27$ [31]),
    .i28(\t/a/regfile/regfile$28$ [31]),
    .i29(\t/a/regfile/regfile$29$ [31]),
    .i3(\t/a/regfile/regfile$3$ [31]),
    .i30(\t/a/regfile/regfile$30$ [31]),
    .i31(\t/a/regfile/regfile$31$ [31]),
    .i4(\t/a/regfile/regfile$4$ [31]),
    .i5(\t/a/regfile/regfile$5$ [31]),
    .i6(\t/a/regfile/regfile$6$ [31]),
    .i7(\t/a/regfile/regfile$7$ [31]),
    .i8(\t/a/regfile/regfile$8$ [31]),
    .i9(\t/a/regfile/regfile$9$ [31]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [31]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b4  (
    .i0(\t/a/regfile/regfile$0$ [4]),
    .i1(\t/a/regfile/regfile$1$ [4]),
    .i10(\t/a/regfile/regfile$10$ [4]),
    .i11(\t/a/regfile/regfile$11$ [4]),
    .i12(\t/a/regfile/regfile$12$ [4]),
    .i13(\t/a/regfile/regfile$13$ [4]),
    .i14(\t/a/regfile/regfile$14$ [4]),
    .i15(\t/a/regfile/regfile$15$ [4]),
    .i16(\t/a/regfile/regfile$16$ [4]),
    .i17(\t/a/regfile/regfile$17$ [4]),
    .i18(\t/a/regfile/regfile$18$ [4]),
    .i19(\t/a/regfile/regfile$19$ [4]),
    .i2(\t/a/regfile/regfile$2$ [4]),
    .i20(\t/a/regfile/regfile$20$ [4]),
    .i21(\t/a/regfile/regfile$21$ [4]),
    .i22(\t/a/regfile/regfile$22$ [4]),
    .i23(\t/a/regfile/regfile$23$ [4]),
    .i24(\t/a/regfile/regfile$24$ [4]),
    .i25(\t/a/regfile/regfile$25$ [4]),
    .i26(\t/a/regfile/regfile$26$ [4]),
    .i27(\t/a/regfile/regfile$27$ [4]),
    .i28(\t/a/regfile/regfile$28$ [4]),
    .i29(\t/a/regfile/regfile$29$ [4]),
    .i3(\t/a/regfile/regfile$3$ [4]),
    .i30(\t/a/regfile/regfile$30$ [4]),
    .i31(\t/a/regfile/regfile$31$ [4]),
    .i4(\t/a/regfile/regfile$4$ [4]),
    .i5(\t/a/regfile/regfile$5$ [4]),
    .i6(\t/a/regfile/regfile$6$ [4]),
    .i7(\t/a/regfile/regfile$7$ [4]),
    .i8(\t/a/regfile/regfile$8$ [4]),
    .i9(\t/a/regfile/regfile$9$ [4]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [4]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b5  (
    .i0(\t/a/regfile/regfile$0$ [5]),
    .i1(\t/a/regfile/regfile$1$ [5]),
    .i10(\t/a/regfile/regfile$10$ [5]),
    .i11(\t/a/regfile/regfile$11$ [5]),
    .i12(\t/a/regfile/regfile$12$ [5]),
    .i13(\t/a/regfile/regfile$13$ [5]),
    .i14(\t/a/regfile/regfile$14$ [5]),
    .i15(\t/a/regfile/regfile$15$ [5]),
    .i16(\t/a/regfile/regfile$16$ [5]),
    .i17(\t/a/regfile/regfile$17$ [5]),
    .i18(\t/a/regfile/regfile$18$ [5]),
    .i19(\t/a/regfile/regfile$19$ [5]),
    .i2(\t/a/regfile/regfile$2$ [5]),
    .i20(\t/a/regfile/regfile$20$ [5]),
    .i21(\t/a/regfile/regfile$21$ [5]),
    .i22(\t/a/regfile/regfile$22$ [5]),
    .i23(\t/a/regfile/regfile$23$ [5]),
    .i24(\t/a/regfile/regfile$24$ [5]),
    .i25(\t/a/regfile/regfile$25$ [5]),
    .i26(\t/a/regfile/regfile$26$ [5]),
    .i27(\t/a/regfile/regfile$27$ [5]),
    .i28(\t/a/regfile/regfile$28$ [5]),
    .i29(\t/a/regfile/regfile$29$ [5]),
    .i3(\t/a/regfile/regfile$3$ [5]),
    .i30(\t/a/regfile/regfile$30$ [5]),
    .i31(\t/a/regfile/regfile$31$ [5]),
    .i4(\t/a/regfile/regfile$4$ [5]),
    .i5(\t/a/regfile/regfile$5$ [5]),
    .i6(\t/a/regfile/regfile$6$ [5]),
    .i7(\t/a/regfile/regfile$7$ [5]),
    .i8(\t/a/regfile/regfile$8$ [5]),
    .i9(\t/a/regfile/regfile$9$ [5]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [5]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b6  (
    .i0(\t/a/regfile/regfile$0$ [6]),
    .i1(\t/a/regfile/regfile$1$ [6]),
    .i10(\t/a/regfile/regfile$10$ [6]),
    .i11(\t/a/regfile/regfile$11$ [6]),
    .i12(\t/a/regfile/regfile$12$ [6]),
    .i13(\t/a/regfile/regfile$13$ [6]),
    .i14(\t/a/regfile/regfile$14$ [6]),
    .i15(\t/a/regfile/regfile$15$ [6]),
    .i16(\t/a/regfile/regfile$16$ [6]),
    .i17(\t/a/regfile/regfile$17$ [6]),
    .i18(\t/a/regfile/regfile$18$ [6]),
    .i19(\t/a/regfile/regfile$19$ [6]),
    .i2(\t/a/regfile/regfile$2$ [6]),
    .i20(\t/a/regfile/regfile$20$ [6]),
    .i21(\t/a/regfile/regfile$21$ [6]),
    .i22(\t/a/regfile/regfile$22$ [6]),
    .i23(\t/a/regfile/regfile$23$ [6]),
    .i24(\t/a/regfile/regfile$24$ [6]),
    .i25(\t/a/regfile/regfile$25$ [6]),
    .i26(\t/a/regfile/regfile$26$ [6]),
    .i27(\t/a/regfile/regfile$27$ [6]),
    .i28(\t/a/regfile/regfile$28$ [6]),
    .i29(\t/a/regfile/regfile$29$ [6]),
    .i3(\t/a/regfile/regfile$3$ [6]),
    .i30(\t/a/regfile/regfile$30$ [6]),
    .i31(\t/a/regfile/regfile$31$ [6]),
    .i4(\t/a/regfile/regfile$4$ [6]),
    .i5(\t/a/regfile/regfile$5$ [6]),
    .i6(\t/a/regfile/regfile$6$ [6]),
    .i7(\t/a/regfile/regfile$7$ [6]),
    .i8(\t/a/regfile/regfile$8$ [6]),
    .i9(\t/a/regfile/regfile$9$ [6]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [6]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b7  (
    .i0(\t/a/regfile/regfile$0$ [7]),
    .i1(\t/a/regfile/regfile$1$ [7]),
    .i10(\t/a/regfile/regfile$10$ [7]),
    .i11(\t/a/regfile/regfile$11$ [7]),
    .i12(\t/a/regfile/regfile$12$ [7]),
    .i13(\t/a/regfile/regfile$13$ [7]),
    .i14(\t/a/regfile/regfile$14$ [7]),
    .i15(\t/a/regfile/regfile$15$ [7]),
    .i16(\t/a/regfile/regfile$16$ [7]),
    .i17(\t/a/regfile/regfile$17$ [7]),
    .i18(\t/a/regfile/regfile$18$ [7]),
    .i19(\t/a/regfile/regfile$19$ [7]),
    .i2(\t/a/regfile/regfile$2$ [7]),
    .i20(\t/a/regfile/regfile$20$ [7]),
    .i21(\t/a/regfile/regfile$21$ [7]),
    .i22(\t/a/regfile/regfile$22$ [7]),
    .i23(\t/a/regfile/regfile$23$ [7]),
    .i24(\t/a/regfile/regfile$24$ [7]),
    .i25(\t/a/regfile/regfile$25$ [7]),
    .i26(\t/a/regfile/regfile$26$ [7]),
    .i27(\t/a/regfile/regfile$27$ [7]),
    .i28(\t/a/regfile/regfile$28$ [7]),
    .i29(\t/a/regfile/regfile$29$ [7]),
    .i3(\t/a/regfile/regfile$3$ [7]),
    .i30(\t/a/regfile/regfile$30$ [7]),
    .i31(\t/a/regfile/regfile$31$ [7]),
    .i4(\t/a/regfile/regfile$4$ [7]),
    .i5(\t/a/regfile/regfile$5$ [7]),
    .i6(\t/a/regfile/regfile$6$ [7]),
    .i7(\t/a/regfile/regfile$7$ [7]),
    .i8(\t/a/regfile/regfile$8$ [7]),
    .i9(\t/a/regfile/regfile$9$ [7]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [7]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b8  (
    .i0(\t/a/regfile/regfile$0$ [8]),
    .i1(\t/a/regfile/regfile$1$ [8]),
    .i10(\t/a/regfile/regfile$10$ [8]),
    .i11(\t/a/regfile/regfile$11$ [8]),
    .i12(\t/a/regfile/regfile$12$ [8]),
    .i13(\t/a/regfile/regfile$13$ [8]),
    .i14(\t/a/regfile/regfile$14$ [8]),
    .i15(\t/a/regfile/regfile$15$ [8]),
    .i16(\t/a/regfile/regfile$16$ [8]),
    .i17(\t/a/regfile/regfile$17$ [8]),
    .i18(\t/a/regfile/regfile$18$ [8]),
    .i19(\t/a/regfile/regfile$19$ [8]),
    .i2(\t/a/regfile/regfile$2$ [8]),
    .i20(\t/a/regfile/regfile$20$ [8]),
    .i21(\t/a/regfile/regfile$21$ [8]),
    .i22(\t/a/regfile/regfile$22$ [8]),
    .i23(\t/a/regfile/regfile$23$ [8]),
    .i24(\t/a/regfile/regfile$24$ [8]),
    .i25(\t/a/regfile/regfile$25$ [8]),
    .i26(\t/a/regfile/regfile$26$ [8]),
    .i27(\t/a/regfile/regfile$27$ [8]),
    .i28(\t/a/regfile/regfile$28$ [8]),
    .i29(\t/a/regfile/regfile$29$ [8]),
    .i3(\t/a/regfile/regfile$3$ [8]),
    .i30(\t/a/regfile/regfile$30$ [8]),
    .i31(\t/a/regfile/regfile$31$ [8]),
    .i4(\t/a/regfile/regfile$4$ [8]),
    .i5(\t/a/regfile/regfile$5$ [8]),
    .i6(\t/a/regfile/regfile$6$ [8]),
    .i7(\t/a/regfile/regfile$7$ [8]),
    .i8(\t/a/regfile/regfile$8$ [8]),
    .i9(\t/a/regfile/regfile$9$ [8]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [8]));  // register.v(16)
  binary_mux_s5_w1 \t/a/regfile/mux0_b9  (
    .i0(\t/a/regfile/regfile$0$ [9]),
    .i1(\t/a/regfile/regfile$1$ [9]),
    .i10(\t/a/regfile/regfile$10$ [9]),
    .i11(\t/a/regfile/regfile$11$ [9]),
    .i12(\t/a/regfile/regfile$12$ [9]),
    .i13(\t/a/regfile/regfile$13$ [9]),
    .i14(\t/a/regfile/regfile$14$ [9]),
    .i15(\t/a/regfile/regfile$15$ [9]),
    .i16(\t/a/regfile/regfile$16$ [9]),
    .i17(\t/a/regfile/regfile$17$ [9]),
    .i18(\t/a/regfile/regfile$18$ [9]),
    .i19(\t/a/regfile/regfile$19$ [9]),
    .i2(\t/a/regfile/regfile$2$ [9]),
    .i20(\t/a/regfile/regfile$20$ [9]),
    .i21(\t/a/regfile/regfile$21$ [9]),
    .i22(\t/a/regfile/regfile$22$ [9]),
    .i23(\t/a/regfile/regfile$23$ [9]),
    .i24(\t/a/regfile/regfile$24$ [9]),
    .i25(\t/a/regfile/regfile$25$ [9]),
    .i26(\t/a/regfile/regfile$26$ [9]),
    .i27(\t/a/regfile/regfile$27$ [9]),
    .i28(\t/a/regfile/regfile$28$ [9]),
    .i29(\t/a/regfile/regfile$29$ [9]),
    .i3(\t/a/regfile/regfile$3$ [9]),
    .i30(\t/a/regfile/regfile$30$ [9]),
    .i31(\t/a/regfile/regfile$31$ [9]),
    .i4(\t/a/regfile/regfile$4$ [9]),
    .i5(\t/a/regfile/regfile$5$ [9]),
    .i6(\t/a/regfile/regfile$6$ [9]),
    .i7(\t/a/regfile/regfile$7$ [9]),
    .i8(\t/a/regfile/regfile$8$ [9]),
    .i9(\t/a/regfile/regfile$9$ [9]),
    .sel(\t/a/ID_rs2 ),
    .o(\t/a/regfile/n5 [9]));  // register.v(16)
  and \t/a/regfile/mux39_b0_sel_is_3  (\t/a/regfile/mux39_b0_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [0]);
  and \t/a/regfile/mux39_b1000_sel_is_3  (\t/a/regfile/mux39_b1000_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [31]);
  and \t/a/regfile/mux39_b100_sel_is_3  (\t/a/regfile/mux39_b100_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [3]);
  and \t/a/regfile/mux39_b128_sel_is_3  (\t/a/regfile/mux39_b128_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [4]);
  and \t/a/regfile/mux39_b160_sel_is_3  (\t/a/regfile/mux39_b160_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [5]);
  and \t/a/regfile/mux39_b192_sel_is_3  (\t/a/regfile/mux39_b192_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [6]);
  and \t/a/regfile/mux39_b224_sel_is_3  (\t/a/regfile/mux39_b224_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [7]);
  and \t/a/regfile/mux39_b256_sel_is_3  (\t/a/regfile/mux39_b256_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [8]);
  and \t/a/regfile/mux39_b288_sel_is_3  (\t/a/regfile/mux39_b288_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [9]);
  and \t/a/regfile/mux39_b320_sel_is_3  (\t/a/regfile/mux39_b320_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [10]);
  and \t/a/regfile/mux39_b32_sel_is_3  (\t/a/regfile/mux39_b32_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [1]);
  and \t/a/regfile/mux39_b352_sel_is_3  (\t/a/regfile/mux39_b352_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [11]);
  and \t/a/regfile/mux39_b384_sel_is_3  (\t/a/regfile/mux39_b384_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [12]);
  and \t/a/regfile/mux39_b416_sel_is_3  (\t/a/regfile/mux39_b416_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [13]);
  and \t/a/regfile/mux39_b448_sel_is_3  (\t/a/regfile/mux39_b448_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [14]);
  and \t/a/regfile/mux39_b480_sel_is_3  (\t/a/regfile/mux39_b480_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [15]);
  and \t/a/regfile/mux39_b512_sel_is_3  (\t/a/regfile/mux39_b512_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [16]);
  and \t/a/regfile/mux39_b544_sel_is_3  (\t/a/regfile/mux39_b544_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [17]);
  and \t/a/regfile/mux39_b576_sel_is_3  (\t/a/regfile/mux39_b576_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [18]);
  and \t/a/regfile/mux39_b608_sel_is_3  (\t/a/regfile/mux39_b608_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [19]);
  and \t/a/regfile/mux39_b640_sel_is_3  (\t/a/regfile/mux39_b640_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [20]);
  and \t/a/regfile/mux39_b64_sel_is_3  (\t/a/regfile/mux39_b64_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [2]);
  and \t/a/regfile/mux39_b672_sel_is_3  (\t/a/regfile/mux39_b672_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [21]);
  and \t/a/regfile/mux39_b704_sel_is_3  (\t/a/regfile/mux39_b704_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [22]);
  and \t/a/regfile/mux39_b736_sel_is_3  (\t/a/regfile/mux39_b736_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [23]);
  and \t/a/regfile/mux39_b768_sel_is_3  (\t/a/regfile/mux39_b768_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [24]);
  and \t/a/regfile/mux39_b800_sel_is_3  (\t/a/regfile/mux39_b800_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [25]);
  and \t/a/regfile/mux39_b832_sel_is_3  (\t/a/regfile/mux39_b832_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [26]);
  and \t/a/regfile/mux39_b864_sel_is_3  (\t/a/regfile/mux39_b864_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [27]);
  and \t/a/regfile/mux39_b896_sel_is_3  (\t/a/regfile/mux39_b896_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [28]);
  and \t/a/regfile/mux39_b928_sel_is_3  (\t/a/regfile/mux39_b928_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [29]);
  and \t/a/regfile/mux39_b960_sel_is_3  (\t/a/regfile/mux39_b960_sel_is_3_o , \t/a/WB_regwritecs , \t/a/regfile/n46 [30]);
  binary_mux_s5_w1 \t/a/regfile/mux40_b0  (
    .i0(\t/a/regfile/regfile$0$ [0]),
    .i1(\t/a/regfile/regfile$1$ [0]),
    .i10(\t/a/regfile/regfile$10$ [0]),
    .i11(\t/a/regfile/regfile$11$ [0]),
    .i12(\t/a/regfile/regfile$12$ [0]),
    .i13(\t/a/regfile/regfile$13$ [0]),
    .i14(\t/a/regfile/regfile$14$ [0]),
    .i15(\t/a/regfile/regfile$15$ [0]),
    .i16(\t/a/regfile/regfile$16$ [0]),
    .i17(\t/a/regfile/regfile$17$ [0]),
    .i18(\t/a/regfile/regfile$18$ [0]),
    .i19(\t/a/regfile/regfile$19$ [0]),
    .i2(\t/a/regfile/regfile$2$ [0]),
    .i20(\t/a/regfile/regfile$20$ [0]),
    .i21(\t/a/regfile/regfile$21$ [0]),
    .i22(\t/a/regfile/regfile$22$ [0]),
    .i23(\t/a/regfile/regfile$23$ [0]),
    .i24(\t/a/regfile/regfile$24$ [0]),
    .i25(\t/a/regfile/regfile$25$ [0]),
    .i26(\t/a/regfile/regfile$26$ [0]),
    .i27(\t/a/regfile/regfile$27$ [0]),
    .i28(\t/a/regfile/regfile$28$ [0]),
    .i29(\t/a/regfile/regfile$29$ [0]),
    .i3(\t/a/regfile/regfile$3$ [0]),
    .i30(\t/a/regfile/regfile$30$ [0]),
    .i31(\t/a/regfile/regfile$31$ [0]),
    .i4(\t/a/regfile/regfile$4$ [0]),
    .i5(\t/a/regfile/regfile$5$ [0]),
    .i6(\t/a/regfile/regfile$6$ [0]),
    .i7(\t/a/regfile/regfile$7$ [0]),
    .i8(\t/a/regfile/regfile$8$ [0]),
    .i9(\t/a/regfile/regfile$9$ [0]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [0]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b1  (
    .i0(\t/a/regfile/regfile$0$ [1]),
    .i1(\t/a/regfile/regfile$1$ [1]),
    .i10(\t/a/regfile/regfile$10$ [1]),
    .i11(\t/a/regfile/regfile$11$ [1]),
    .i12(\t/a/regfile/regfile$12$ [1]),
    .i13(\t/a/regfile/regfile$13$ [1]),
    .i14(\t/a/regfile/regfile$14$ [1]),
    .i15(\t/a/regfile/regfile$15$ [1]),
    .i16(\t/a/regfile/regfile$16$ [1]),
    .i17(\t/a/regfile/regfile$17$ [1]),
    .i18(\t/a/regfile/regfile$18$ [1]),
    .i19(\t/a/regfile/regfile$19$ [1]),
    .i2(\t/a/regfile/regfile$2$ [1]),
    .i20(\t/a/regfile/regfile$20$ [1]),
    .i21(\t/a/regfile/regfile$21$ [1]),
    .i22(\t/a/regfile/regfile$22$ [1]),
    .i23(\t/a/regfile/regfile$23$ [1]),
    .i24(\t/a/regfile/regfile$24$ [1]),
    .i25(\t/a/regfile/regfile$25$ [1]),
    .i26(\t/a/regfile/regfile$26$ [1]),
    .i27(\t/a/regfile/regfile$27$ [1]),
    .i28(\t/a/regfile/regfile$28$ [1]),
    .i29(\t/a/regfile/regfile$29$ [1]),
    .i3(\t/a/regfile/regfile$3$ [1]),
    .i30(\t/a/regfile/regfile$30$ [1]),
    .i31(\t/a/regfile/regfile$31$ [1]),
    .i4(\t/a/regfile/regfile$4$ [1]),
    .i5(\t/a/regfile/regfile$5$ [1]),
    .i6(\t/a/regfile/regfile$6$ [1]),
    .i7(\t/a/regfile/regfile$7$ [1]),
    .i8(\t/a/regfile/regfile$8$ [1]),
    .i9(\t/a/regfile/regfile$9$ [1]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [1]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b10  (
    .i0(\t/a/regfile/regfile$0$ [10]),
    .i1(\t/a/regfile/regfile$1$ [10]),
    .i10(\t/a/regfile/regfile$10$ [10]),
    .i11(\t/a/regfile/regfile$11$ [10]),
    .i12(\t/a/regfile/regfile$12$ [10]),
    .i13(\t/a/regfile/regfile$13$ [10]),
    .i14(\t/a/regfile/regfile$14$ [10]),
    .i15(\t/a/regfile/regfile$15$ [10]),
    .i16(\t/a/regfile/regfile$16$ [10]),
    .i17(\t/a/regfile/regfile$17$ [10]),
    .i18(\t/a/regfile/regfile$18$ [10]),
    .i19(\t/a/regfile/regfile$19$ [10]),
    .i2(\t/a/regfile/regfile$2$ [10]),
    .i20(\t/a/regfile/regfile$20$ [10]),
    .i21(\t/a/regfile/regfile$21$ [10]),
    .i22(\t/a/regfile/regfile$22$ [10]),
    .i23(\t/a/regfile/regfile$23$ [10]),
    .i24(\t/a/regfile/regfile$24$ [10]),
    .i25(\t/a/regfile/regfile$25$ [10]),
    .i26(\t/a/regfile/regfile$26$ [10]),
    .i27(\t/a/regfile/regfile$27$ [10]),
    .i28(\t/a/regfile/regfile$28$ [10]),
    .i29(\t/a/regfile/regfile$29$ [10]),
    .i3(\t/a/regfile/regfile$3$ [10]),
    .i30(\t/a/regfile/regfile$30$ [10]),
    .i31(\t/a/regfile/regfile$31$ [10]),
    .i4(\t/a/regfile/regfile$4$ [10]),
    .i5(\t/a/regfile/regfile$5$ [10]),
    .i6(\t/a/regfile/regfile$6$ [10]),
    .i7(\t/a/regfile/regfile$7$ [10]),
    .i8(\t/a/regfile/regfile$8$ [10]),
    .i9(\t/a/regfile/regfile$9$ [10]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [10]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b11  (
    .i0(\t/a/regfile/regfile$0$ [11]),
    .i1(\t/a/regfile/regfile$1$ [11]),
    .i10(\t/a/regfile/regfile$10$ [11]),
    .i11(\t/a/regfile/regfile$11$ [11]),
    .i12(\t/a/regfile/regfile$12$ [11]),
    .i13(\t/a/regfile/regfile$13$ [11]),
    .i14(\t/a/regfile/regfile$14$ [11]),
    .i15(\t/a/regfile/regfile$15$ [11]),
    .i16(\t/a/regfile/regfile$16$ [11]),
    .i17(\t/a/regfile/regfile$17$ [11]),
    .i18(\t/a/regfile/regfile$18$ [11]),
    .i19(\t/a/regfile/regfile$19$ [11]),
    .i2(\t/a/regfile/regfile$2$ [11]),
    .i20(\t/a/regfile/regfile$20$ [11]),
    .i21(\t/a/regfile/regfile$21$ [11]),
    .i22(\t/a/regfile/regfile$22$ [11]),
    .i23(\t/a/regfile/regfile$23$ [11]),
    .i24(\t/a/regfile/regfile$24$ [11]),
    .i25(\t/a/regfile/regfile$25$ [11]),
    .i26(\t/a/regfile/regfile$26$ [11]),
    .i27(\t/a/regfile/regfile$27$ [11]),
    .i28(\t/a/regfile/regfile$28$ [11]),
    .i29(\t/a/regfile/regfile$29$ [11]),
    .i3(\t/a/regfile/regfile$3$ [11]),
    .i30(\t/a/regfile/regfile$30$ [11]),
    .i31(\t/a/regfile/regfile$31$ [11]),
    .i4(\t/a/regfile/regfile$4$ [11]),
    .i5(\t/a/regfile/regfile$5$ [11]),
    .i6(\t/a/regfile/regfile$6$ [11]),
    .i7(\t/a/regfile/regfile$7$ [11]),
    .i8(\t/a/regfile/regfile$8$ [11]),
    .i9(\t/a/regfile/regfile$9$ [11]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [11]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b12  (
    .i0(\t/a/regfile/regfile$0$ [12]),
    .i1(\t/a/regfile/regfile$1$ [12]),
    .i10(\t/a/regfile/regfile$10$ [12]),
    .i11(\t/a/regfile/regfile$11$ [12]),
    .i12(\t/a/regfile/regfile$12$ [12]),
    .i13(\t/a/regfile/regfile$13$ [12]),
    .i14(\t/a/regfile/regfile$14$ [12]),
    .i15(\t/a/regfile/regfile$15$ [12]),
    .i16(\t/a/regfile/regfile$16$ [12]),
    .i17(\t/a/regfile/regfile$17$ [12]),
    .i18(\t/a/regfile/regfile$18$ [12]),
    .i19(\t/a/regfile/regfile$19$ [12]),
    .i2(\t/a/regfile/regfile$2$ [12]),
    .i20(\t/a/regfile/regfile$20$ [12]),
    .i21(\t/a/regfile/regfile$21$ [12]),
    .i22(\t/a/regfile/regfile$22$ [12]),
    .i23(\t/a/regfile/regfile$23$ [12]),
    .i24(\t/a/regfile/regfile$24$ [12]),
    .i25(\t/a/regfile/regfile$25$ [12]),
    .i26(\t/a/regfile/regfile$26$ [12]),
    .i27(\t/a/regfile/regfile$27$ [12]),
    .i28(\t/a/regfile/regfile$28$ [12]),
    .i29(\t/a/regfile/regfile$29$ [12]),
    .i3(\t/a/regfile/regfile$3$ [12]),
    .i30(\t/a/regfile/regfile$30$ [12]),
    .i31(\t/a/regfile/regfile$31$ [12]),
    .i4(\t/a/regfile/regfile$4$ [12]),
    .i5(\t/a/regfile/regfile$5$ [12]),
    .i6(\t/a/regfile/regfile$6$ [12]),
    .i7(\t/a/regfile/regfile$7$ [12]),
    .i8(\t/a/regfile/regfile$8$ [12]),
    .i9(\t/a/regfile/regfile$9$ [12]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [12]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b13  (
    .i0(\t/a/regfile/regfile$0$ [13]),
    .i1(\t/a/regfile/regfile$1$ [13]),
    .i10(\t/a/regfile/regfile$10$ [13]),
    .i11(\t/a/regfile/regfile$11$ [13]),
    .i12(\t/a/regfile/regfile$12$ [13]),
    .i13(\t/a/regfile/regfile$13$ [13]),
    .i14(\t/a/regfile/regfile$14$ [13]),
    .i15(\t/a/regfile/regfile$15$ [13]),
    .i16(\t/a/regfile/regfile$16$ [13]),
    .i17(\t/a/regfile/regfile$17$ [13]),
    .i18(\t/a/regfile/regfile$18$ [13]),
    .i19(\t/a/regfile/regfile$19$ [13]),
    .i2(\t/a/regfile/regfile$2$ [13]),
    .i20(\t/a/regfile/regfile$20$ [13]),
    .i21(\t/a/regfile/regfile$21$ [13]),
    .i22(\t/a/regfile/regfile$22$ [13]),
    .i23(\t/a/regfile/regfile$23$ [13]),
    .i24(\t/a/regfile/regfile$24$ [13]),
    .i25(\t/a/regfile/regfile$25$ [13]),
    .i26(\t/a/regfile/regfile$26$ [13]),
    .i27(\t/a/regfile/regfile$27$ [13]),
    .i28(\t/a/regfile/regfile$28$ [13]),
    .i29(\t/a/regfile/regfile$29$ [13]),
    .i3(\t/a/regfile/regfile$3$ [13]),
    .i30(\t/a/regfile/regfile$30$ [13]),
    .i31(\t/a/regfile/regfile$31$ [13]),
    .i4(\t/a/regfile/regfile$4$ [13]),
    .i5(\t/a/regfile/regfile$5$ [13]),
    .i6(\t/a/regfile/regfile$6$ [13]),
    .i7(\t/a/regfile/regfile$7$ [13]),
    .i8(\t/a/regfile/regfile$8$ [13]),
    .i9(\t/a/regfile/regfile$9$ [13]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [13]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b14  (
    .i0(\t/a/regfile/regfile$0$ [14]),
    .i1(\t/a/regfile/regfile$1$ [14]),
    .i10(\t/a/regfile/regfile$10$ [14]),
    .i11(\t/a/regfile/regfile$11$ [14]),
    .i12(\t/a/regfile/regfile$12$ [14]),
    .i13(\t/a/regfile/regfile$13$ [14]),
    .i14(\t/a/regfile/regfile$14$ [14]),
    .i15(\t/a/regfile/regfile$15$ [14]),
    .i16(\t/a/regfile/regfile$16$ [14]),
    .i17(\t/a/regfile/regfile$17$ [14]),
    .i18(\t/a/regfile/regfile$18$ [14]),
    .i19(\t/a/regfile/regfile$19$ [14]),
    .i2(\t/a/regfile/regfile$2$ [14]),
    .i20(\t/a/regfile/regfile$20$ [14]),
    .i21(\t/a/regfile/regfile$21$ [14]),
    .i22(\t/a/regfile/regfile$22$ [14]),
    .i23(\t/a/regfile/regfile$23$ [14]),
    .i24(\t/a/regfile/regfile$24$ [14]),
    .i25(\t/a/regfile/regfile$25$ [14]),
    .i26(\t/a/regfile/regfile$26$ [14]),
    .i27(\t/a/regfile/regfile$27$ [14]),
    .i28(\t/a/regfile/regfile$28$ [14]),
    .i29(\t/a/regfile/regfile$29$ [14]),
    .i3(\t/a/regfile/regfile$3$ [14]),
    .i30(\t/a/regfile/regfile$30$ [14]),
    .i31(\t/a/regfile/regfile$31$ [14]),
    .i4(\t/a/regfile/regfile$4$ [14]),
    .i5(\t/a/regfile/regfile$5$ [14]),
    .i6(\t/a/regfile/regfile$6$ [14]),
    .i7(\t/a/regfile/regfile$7$ [14]),
    .i8(\t/a/regfile/regfile$8$ [14]),
    .i9(\t/a/regfile/regfile$9$ [14]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [14]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b15  (
    .i0(\t/a/regfile/regfile$0$ [15]),
    .i1(\t/a/regfile/regfile$1$ [15]),
    .i10(\t/a/regfile/regfile$10$ [15]),
    .i11(\t/a/regfile/regfile$11$ [15]),
    .i12(\t/a/regfile/regfile$12$ [15]),
    .i13(\t/a/regfile/regfile$13$ [15]),
    .i14(\t/a/regfile/regfile$14$ [15]),
    .i15(\t/a/regfile/regfile$15$ [15]),
    .i16(\t/a/regfile/regfile$16$ [15]),
    .i17(\t/a/regfile/regfile$17$ [15]),
    .i18(\t/a/regfile/regfile$18$ [15]),
    .i19(\t/a/regfile/regfile$19$ [15]),
    .i2(\t/a/regfile/regfile$2$ [15]),
    .i20(\t/a/regfile/regfile$20$ [15]),
    .i21(\t/a/regfile/regfile$21$ [15]),
    .i22(\t/a/regfile/regfile$22$ [15]),
    .i23(\t/a/regfile/regfile$23$ [15]),
    .i24(\t/a/regfile/regfile$24$ [15]),
    .i25(\t/a/regfile/regfile$25$ [15]),
    .i26(\t/a/regfile/regfile$26$ [15]),
    .i27(\t/a/regfile/regfile$27$ [15]),
    .i28(\t/a/regfile/regfile$28$ [15]),
    .i29(\t/a/regfile/regfile$29$ [15]),
    .i3(\t/a/regfile/regfile$3$ [15]),
    .i30(\t/a/regfile/regfile$30$ [15]),
    .i31(\t/a/regfile/regfile$31$ [15]),
    .i4(\t/a/regfile/regfile$4$ [15]),
    .i5(\t/a/regfile/regfile$5$ [15]),
    .i6(\t/a/regfile/regfile$6$ [15]),
    .i7(\t/a/regfile/regfile$7$ [15]),
    .i8(\t/a/regfile/regfile$8$ [15]),
    .i9(\t/a/regfile/regfile$9$ [15]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [15]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b16  (
    .i0(\t/a/regfile/regfile$0$ [16]),
    .i1(\t/a/regfile/regfile$1$ [16]),
    .i10(\t/a/regfile/regfile$10$ [16]),
    .i11(\t/a/regfile/regfile$11$ [16]),
    .i12(\t/a/regfile/regfile$12$ [16]),
    .i13(\t/a/regfile/regfile$13$ [16]),
    .i14(\t/a/regfile/regfile$14$ [16]),
    .i15(\t/a/regfile/regfile$15$ [16]),
    .i16(\t/a/regfile/regfile$16$ [16]),
    .i17(\t/a/regfile/regfile$17$ [16]),
    .i18(\t/a/regfile/regfile$18$ [16]),
    .i19(\t/a/regfile/regfile$19$ [16]),
    .i2(\t/a/regfile/regfile$2$ [16]),
    .i20(\t/a/regfile/regfile$20$ [16]),
    .i21(\t/a/regfile/regfile$21$ [16]),
    .i22(\t/a/regfile/regfile$22$ [16]),
    .i23(\t/a/regfile/regfile$23$ [16]),
    .i24(\t/a/regfile/regfile$24$ [16]),
    .i25(\t/a/regfile/regfile$25$ [16]),
    .i26(\t/a/regfile/regfile$26$ [16]),
    .i27(\t/a/regfile/regfile$27$ [16]),
    .i28(\t/a/regfile/regfile$28$ [16]),
    .i29(\t/a/regfile/regfile$29$ [16]),
    .i3(\t/a/regfile/regfile$3$ [16]),
    .i30(\t/a/regfile/regfile$30$ [16]),
    .i31(\t/a/regfile/regfile$31$ [16]),
    .i4(\t/a/regfile/regfile$4$ [16]),
    .i5(\t/a/regfile/regfile$5$ [16]),
    .i6(\t/a/regfile/regfile$6$ [16]),
    .i7(\t/a/regfile/regfile$7$ [16]),
    .i8(\t/a/regfile/regfile$8$ [16]),
    .i9(\t/a/regfile/regfile$9$ [16]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [16]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b17  (
    .i0(\t/a/regfile/regfile$0$ [17]),
    .i1(\t/a/regfile/regfile$1$ [17]),
    .i10(\t/a/regfile/regfile$10$ [17]),
    .i11(\t/a/regfile/regfile$11$ [17]),
    .i12(\t/a/regfile/regfile$12$ [17]),
    .i13(\t/a/regfile/regfile$13$ [17]),
    .i14(\t/a/regfile/regfile$14$ [17]),
    .i15(\t/a/regfile/regfile$15$ [17]),
    .i16(\t/a/regfile/regfile$16$ [17]),
    .i17(\t/a/regfile/regfile$17$ [17]),
    .i18(\t/a/regfile/regfile$18$ [17]),
    .i19(\t/a/regfile/regfile$19$ [17]),
    .i2(\t/a/regfile/regfile$2$ [17]),
    .i20(\t/a/regfile/regfile$20$ [17]),
    .i21(\t/a/regfile/regfile$21$ [17]),
    .i22(\t/a/regfile/regfile$22$ [17]),
    .i23(\t/a/regfile/regfile$23$ [17]),
    .i24(\t/a/regfile/regfile$24$ [17]),
    .i25(\t/a/regfile/regfile$25$ [17]),
    .i26(\t/a/regfile/regfile$26$ [17]),
    .i27(\t/a/regfile/regfile$27$ [17]),
    .i28(\t/a/regfile/regfile$28$ [17]),
    .i29(\t/a/regfile/regfile$29$ [17]),
    .i3(\t/a/regfile/regfile$3$ [17]),
    .i30(\t/a/regfile/regfile$30$ [17]),
    .i31(\t/a/regfile/regfile$31$ [17]),
    .i4(\t/a/regfile/regfile$4$ [17]),
    .i5(\t/a/regfile/regfile$5$ [17]),
    .i6(\t/a/regfile/regfile$6$ [17]),
    .i7(\t/a/regfile/regfile$7$ [17]),
    .i8(\t/a/regfile/regfile$8$ [17]),
    .i9(\t/a/regfile/regfile$9$ [17]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [17]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b18  (
    .i0(\t/a/regfile/regfile$0$ [18]),
    .i1(\t/a/regfile/regfile$1$ [18]),
    .i10(\t/a/regfile/regfile$10$ [18]),
    .i11(\t/a/regfile/regfile$11$ [18]),
    .i12(\t/a/regfile/regfile$12$ [18]),
    .i13(\t/a/regfile/regfile$13$ [18]),
    .i14(\t/a/regfile/regfile$14$ [18]),
    .i15(\t/a/regfile/regfile$15$ [18]),
    .i16(\t/a/regfile/regfile$16$ [18]),
    .i17(\t/a/regfile/regfile$17$ [18]),
    .i18(\t/a/regfile/regfile$18$ [18]),
    .i19(\t/a/regfile/regfile$19$ [18]),
    .i2(\t/a/regfile/regfile$2$ [18]),
    .i20(\t/a/regfile/regfile$20$ [18]),
    .i21(\t/a/regfile/regfile$21$ [18]),
    .i22(\t/a/regfile/regfile$22$ [18]),
    .i23(\t/a/regfile/regfile$23$ [18]),
    .i24(\t/a/regfile/regfile$24$ [18]),
    .i25(\t/a/regfile/regfile$25$ [18]),
    .i26(\t/a/regfile/regfile$26$ [18]),
    .i27(\t/a/regfile/regfile$27$ [18]),
    .i28(\t/a/regfile/regfile$28$ [18]),
    .i29(\t/a/regfile/regfile$29$ [18]),
    .i3(\t/a/regfile/regfile$3$ [18]),
    .i30(\t/a/regfile/regfile$30$ [18]),
    .i31(\t/a/regfile/regfile$31$ [18]),
    .i4(\t/a/regfile/regfile$4$ [18]),
    .i5(\t/a/regfile/regfile$5$ [18]),
    .i6(\t/a/regfile/regfile$6$ [18]),
    .i7(\t/a/regfile/regfile$7$ [18]),
    .i8(\t/a/regfile/regfile$8$ [18]),
    .i9(\t/a/regfile/regfile$9$ [18]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [18]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b19  (
    .i0(\t/a/regfile/regfile$0$ [19]),
    .i1(\t/a/regfile/regfile$1$ [19]),
    .i10(\t/a/regfile/regfile$10$ [19]),
    .i11(\t/a/regfile/regfile$11$ [19]),
    .i12(\t/a/regfile/regfile$12$ [19]),
    .i13(\t/a/regfile/regfile$13$ [19]),
    .i14(\t/a/regfile/regfile$14$ [19]),
    .i15(\t/a/regfile/regfile$15$ [19]),
    .i16(\t/a/regfile/regfile$16$ [19]),
    .i17(\t/a/regfile/regfile$17$ [19]),
    .i18(\t/a/regfile/regfile$18$ [19]),
    .i19(\t/a/regfile/regfile$19$ [19]),
    .i2(\t/a/regfile/regfile$2$ [19]),
    .i20(\t/a/regfile/regfile$20$ [19]),
    .i21(\t/a/regfile/regfile$21$ [19]),
    .i22(\t/a/regfile/regfile$22$ [19]),
    .i23(\t/a/regfile/regfile$23$ [19]),
    .i24(\t/a/regfile/regfile$24$ [19]),
    .i25(\t/a/regfile/regfile$25$ [19]),
    .i26(\t/a/regfile/regfile$26$ [19]),
    .i27(\t/a/regfile/regfile$27$ [19]),
    .i28(\t/a/regfile/regfile$28$ [19]),
    .i29(\t/a/regfile/regfile$29$ [19]),
    .i3(\t/a/regfile/regfile$3$ [19]),
    .i30(\t/a/regfile/regfile$30$ [19]),
    .i31(\t/a/regfile/regfile$31$ [19]),
    .i4(\t/a/regfile/regfile$4$ [19]),
    .i5(\t/a/regfile/regfile$5$ [19]),
    .i6(\t/a/regfile/regfile$6$ [19]),
    .i7(\t/a/regfile/regfile$7$ [19]),
    .i8(\t/a/regfile/regfile$8$ [19]),
    .i9(\t/a/regfile/regfile$9$ [19]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [19]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b2  (
    .i0(\t/a/regfile/regfile$0$ [2]),
    .i1(\t/a/regfile/regfile$1$ [2]),
    .i10(\t/a/regfile/regfile$10$ [2]),
    .i11(\t/a/regfile/regfile$11$ [2]),
    .i12(\t/a/regfile/regfile$12$ [2]),
    .i13(\t/a/regfile/regfile$13$ [2]),
    .i14(\t/a/regfile/regfile$14$ [2]),
    .i15(\t/a/regfile/regfile$15$ [2]),
    .i16(\t/a/regfile/regfile$16$ [2]),
    .i17(\t/a/regfile/regfile$17$ [2]),
    .i18(\t/a/regfile/regfile$18$ [2]),
    .i19(\t/a/regfile/regfile$19$ [2]),
    .i2(\t/a/regfile/regfile$2$ [2]),
    .i20(\t/a/regfile/regfile$20$ [2]),
    .i21(\t/a/regfile/regfile$21$ [2]),
    .i22(\t/a/regfile/regfile$22$ [2]),
    .i23(\t/a/regfile/regfile$23$ [2]),
    .i24(\t/a/regfile/regfile$24$ [2]),
    .i25(\t/a/regfile/regfile$25$ [2]),
    .i26(\t/a/regfile/regfile$26$ [2]),
    .i27(\t/a/regfile/regfile$27$ [2]),
    .i28(\t/a/regfile/regfile$28$ [2]),
    .i29(\t/a/regfile/regfile$29$ [2]),
    .i3(\t/a/regfile/regfile$3$ [2]),
    .i30(\t/a/regfile/regfile$30$ [2]),
    .i31(\t/a/regfile/regfile$31$ [2]),
    .i4(\t/a/regfile/regfile$4$ [2]),
    .i5(\t/a/regfile/regfile$5$ [2]),
    .i6(\t/a/regfile/regfile$6$ [2]),
    .i7(\t/a/regfile/regfile$7$ [2]),
    .i8(\t/a/regfile/regfile$8$ [2]),
    .i9(\t/a/regfile/regfile$9$ [2]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [2]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b20  (
    .i0(\t/a/regfile/regfile$0$ [20]),
    .i1(\t/a/regfile/regfile$1$ [20]),
    .i10(\t/a/regfile/regfile$10$ [20]),
    .i11(\t/a/regfile/regfile$11$ [20]),
    .i12(\t/a/regfile/regfile$12$ [20]),
    .i13(\t/a/regfile/regfile$13$ [20]),
    .i14(\t/a/regfile/regfile$14$ [20]),
    .i15(\t/a/regfile/regfile$15$ [20]),
    .i16(\t/a/regfile/regfile$16$ [20]),
    .i17(\t/a/regfile/regfile$17$ [20]),
    .i18(\t/a/regfile/regfile$18$ [20]),
    .i19(\t/a/regfile/regfile$19$ [20]),
    .i2(\t/a/regfile/regfile$2$ [20]),
    .i20(\t/a/regfile/regfile$20$ [20]),
    .i21(\t/a/regfile/regfile$21$ [20]),
    .i22(\t/a/regfile/regfile$22$ [20]),
    .i23(\t/a/regfile/regfile$23$ [20]),
    .i24(\t/a/regfile/regfile$24$ [20]),
    .i25(\t/a/regfile/regfile$25$ [20]),
    .i26(\t/a/regfile/regfile$26$ [20]),
    .i27(\t/a/regfile/regfile$27$ [20]),
    .i28(\t/a/regfile/regfile$28$ [20]),
    .i29(\t/a/regfile/regfile$29$ [20]),
    .i3(\t/a/regfile/regfile$3$ [20]),
    .i30(\t/a/regfile/regfile$30$ [20]),
    .i31(\t/a/regfile/regfile$31$ [20]),
    .i4(\t/a/regfile/regfile$4$ [20]),
    .i5(\t/a/regfile/regfile$5$ [20]),
    .i6(\t/a/regfile/regfile$6$ [20]),
    .i7(\t/a/regfile/regfile$7$ [20]),
    .i8(\t/a/regfile/regfile$8$ [20]),
    .i9(\t/a/regfile/regfile$9$ [20]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [20]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b21  (
    .i0(\t/a/regfile/regfile$0$ [21]),
    .i1(\t/a/regfile/regfile$1$ [21]),
    .i10(\t/a/regfile/regfile$10$ [21]),
    .i11(\t/a/regfile/regfile$11$ [21]),
    .i12(\t/a/regfile/regfile$12$ [21]),
    .i13(\t/a/regfile/regfile$13$ [21]),
    .i14(\t/a/regfile/regfile$14$ [21]),
    .i15(\t/a/regfile/regfile$15$ [21]),
    .i16(\t/a/regfile/regfile$16$ [21]),
    .i17(\t/a/regfile/regfile$17$ [21]),
    .i18(\t/a/regfile/regfile$18$ [21]),
    .i19(\t/a/regfile/regfile$19$ [21]),
    .i2(\t/a/regfile/regfile$2$ [21]),
    .i20(\t/a/regfile/regfile$20$ [21]),
    .i21(\t/a/regfile/regfile$21$ [21]),
    .i22(\t/a/regfile/regfile$22$ [21]),
    .i23(\t/a/regfile/regfile$23$ [21]),
    .i24(\t/a/regfile/regfile$24$ [21]),
    .i25(\t/a/regfile/regfile$25$ [21]),
    .i26(\t/a/regfile/regfile$26$ [21]),
    .i27(\t/a/regfile/regfile$27$ [21]),
    .i28(\t/a/regfile/regfile$28$ [21]),
    .i29(\t/a/regfile/regfile$29$ [21]),
    .i3(\t/a/regfile/regfile$3$ [21]),
    .i30(\t/a/regfile/regfile$30$ [21]),
    .i31(\t/a/regfile/regfile$31$ [21]),
    .i4(\t/a/regfile/regfile$4$ [21]),
    .i5(\t/a/regfile/regfile$5$ [21]),
    .i6(\t/a/regfile/regfile$6$ [21]),
    .i7(\t/a/regfile/regfile$7$ [21]),
    .i8(\t/a/regfile/regfile$8$ [21]),
    .i9(\t/a/regfile/regfile$9$ [21]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [21]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b22  (
    .i0(\t/a/regfile/regfile$0$ [22]),
    .i1(\t/a/regfile/regfile$1$ [22]),
    .i10(\t/a/regfile/regfile$10$ [22]),
    .i11(\t/a/regfile/regfile$11$ [22]),
    .i12(\t/a/regfile/regfile$12$ [22]),
    .i13(\t/a/regfile/regfile$13$ [22]),
    .i14(\t/a/regfile/regfile$14$ [22]),
    .i15(\t/a/regfile/regfile$15$ [22]),
    .i16(\t/a/regfile/regfile$16$ [22]),
    .i17(\t/a/regfile/regfile$17$ [22]),
    .i18(\t/a/regfile/regfile$18$ [22]),
    .i19(\t/a/regfile/regfile$19$ [22]),
    .i2(\t/a/regfile/regfile$2$ [22]),
    .i20(\t/a/regfile/regfile$20$ [22]),
    .i21(\t/a/regfile/regfile$21$ [22]),
    .i22(\t/a/regfile/regfile$22$ [22]),
    .i23(\t/a/regfile/regfile$23$ [22]),
    .i24(\t/a/regfile/regfile$24$ [22]),
    .i25(\t/a/regfile/regfile$25$ [22]),
    .i26(\t/a/regfile/regfile$26$ [22]),
    .i27(\t/a/regfile/regfile$27$ [22]),
    .i28(\t/a/regfile/regfile$28$ [22]),
    .i29(\t/a/regfile/regfile$29$ [22]),
    .i3(\t/a/regfile/regfile$3$ [22]),
    .i30(\t/a/regfile/regfile$30$ [22]),
    .i31(\t/a/regfile/regfile$31$ [22]),
    .i4(\t/a/regfile/regfile$4$ [22]),
    .i5(\t/a/regfile/regfile$5$ [22]),
    .i6(\t/a/regfile/regfile$6$ [22]),
    .i7(\t/a/regfile/regfile$7$ [22]),
    .i8(\t/a/regfile/regfile$8$ [22]),
    .i9(\t/a/regfile/regfile$9$ [22]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [22]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b23  (
    .i0(\t/a/regfile/regfile$0$ [23]),
    .i1(\t/a/regfile/regfile$1$ [23]),
    .i10(\t/a/regfile/regfile$10$ [23]),
    .i11(\t/a/regfile/regfile$11$ [23]),
    .i12(\t/a/regfile/regfile$12$ [23]),
    .i13(\t/a/regfile/regfile$13$ [23]),
    .i14(\t/a/regfile/regfile$14$ [23]),
    .i15(\t/a/regfile/regfile$15$ [23]),
    .i16(\t/a/regfile/regfile$16$ [23]),
    .i17(\t/a/regfile/regfile$17$ [23]),
    .i18(\t/a/regfile/regfile$18$ [23]),
    .i19(\t/a/regfile/regfile$19$ [23]),
    .i2(\t/a/regfile/regfile$2$ [23]),
    .i20(\t/a/regfile/regfile$20$ [23]),
    .i21(\t/a/regfile/regfile$21$ [23]),
    .i22(\t/a/regfile/regfile$22$ [23]),
    .i23(\t/a/regfile/regfile$23$ [23]),
    .i24(\t/a/regfile/regfile$24$ [23]),
    .i25(\t/a/regfile/regfile$25$ [23]),
    .i26(\t/a/regfile/regfile$26$ [23]),
    .i27(\t/a/regfile/regfile$27$ [23]),
    .i28(\t/a/regfile/regfile$28$ [23]),
    .i29(\t/a/regfile/regfile$29$ [23]),
    .i3(\t/a/regfile/regfile$3$ [23]),
    .i30(\t/a/regfile/regfile$30$ [23]),
    .i31(\t/a/regfile/regfile$31$ [23]),
    .i4(\t/a/regfile/regfile$4$ [23]),
    .i5(\t/a/regfile/regfile$5$ [23]),
    .i6(\t/a/regfile/regfile$6$ [23]),
    .i7(\t/a/regfile/regfile$7$ [23]),
    .i8(\t/a/regfile/regfile$8$ [23]),
    .i9(\t/a/regfile/regfile$9$ [23]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [23]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b24  (
    .i0(\t/a/regfile/regfile$0$ [24]),
    .i1(\t/a/regfile/regfile$1$ [24]),
    .i10(\t/a/regfile/regfile$10$ [24]),
    .i11(\t/a/regfile/regfile$11$ [24]),
    .i12(\t/a/regfile/regfile$12$ [24]),
    .i13(\t/a/regfile/regfile$13$ [24]),
    .i14(\t/a/regfile/regfile$14$ [24]),
    .i15(\t/a/regfile/regfile$15$ [24]),
    .i16(\t/a/regfile/regfile$16$ [24]),
    .i17(\t/a/regfile/regfile$17$ [24]),
    .i18(\t/a/regfile/regfile$18$ [24]),
    .i19(\t/a/regfile/regfile$19$ [24]),
    .i2(\t/a/regfile/regfile$2$ [24]),
    .i20(\t/a/regfile/regfile$20$ [24]),
    .i21(\t/a/regfile/regfile$21$ [24]),
    .i22(\t/a/regfile/regfile$22$ [24]),
    .i23(\t/a/regfile/regfile$23$ [24]),
    .i24(\t/a/regfile/regfile$24$ [24]),
    .i25(\t/a/regfile/regfile$25$ [24]),
    .i26(\t/a/regfile/regfile$26$ [24]),
    .i27(\t/a/regfile/regfile$27$ [24]),
    .i28(\t/a/regfile/regfile$28$ [24]),
    .i29(\t/a/regfile/regfile$29$ [24]),
    .i3(\t/a/regfile/regfile$3$ [24]),
    .i30(\t/a/regfile/regfile$30$ [24]),
    .i31(\t/a/regfile/regfile$31$ [24]),
    .i4(\t/a/regfile/regfile$4$ [24]),
    .i5(\t/a/regfile/regfile$5$ [24]),
    .i6(\t/a/regfile/regfile$6$ [24]),
    .i7(\t/a/regfile/regfile$7$ [24]),
    .i8(\t/a/regfile/regfile$8$ [24]),
    .i9(\t/a/regfile/regfile$9$ [24]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [24]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b25  (
    .i0(\t/a/regfile/regfile$0$ [25]),
    .i1(\t/a/regfile/regfile$1$ [25]),
    .i10(\t/a/regfile/regfile$10$ [25]),
    .i11(\t/a/regfile/regfile$11$ [25]),
    .i12(\t/a/regfile/regfile$12$ [25]),
    .i13(\t/a/regfile/regfile$13$ [25]),
    .i14(\t/a/regfile/regfile$14$ [25]),
    .i15(\t/a/regfile/regfile$15$ [25]),
    .i16(\t/a/regfile/regfile$16$ [25]),
    .i17(\t/a/regfile/regfile$17$ [25]),
    .i18(\t/a/regfile/regfile$18$ [25]),
    .i19(\t/a/regfile/regfile$19$ [25]),
    .i2(\t/a/regfile/regfile$2$ [25]),
    .i20(\t/a/regfile/regfile$20$ [25]),
    .i21(\t/a/regfile/regfile$21$ [25]),
    .i22(\t/a/regfile/regfile$22$ [25]),
    .i23(\t/a/regfile/regfile$23$ [25]),
    .i24(\t/a/regfile/regfile$24$ [25]),
    .i25(\t/a/regfile/regfile$25$ [25]),
    .i26(\t/a/regfile/regfile$26$ [25]),
    .i27(\t/a/regfile/regfile$27$ [25]),
    .i28(\t/a/regfile/regfile$28$ [25]),
    .i29(\t/a/regfile/regfile$29$ [25]),
    .i3(\t/a/regfile/regfile$3$ [25]),
    .i30(\t/a/regfile/regfile$30$ [25]),
    .i31(\t/a/regfile/regfile$31$ [25]),
    .i4(\t/a/regfile/regfile$4$ [25]),
    .i5(\t/a/regfile/regfile$5$ [25]),
    .i6(\t/a/regfile/regfile$6$ [25]),
    .i7(\t/a/regfile/regfile$7$ [25]),
    .i8(\t/a/regfile/regfile$8$ [25]),
    .i9(\t/a/regfile/regfile$9$ [25]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [25]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b26  (
    .i0(\t/a/regfile/regfile$0$ [26]),
    .i1(\t/a/regfile/regfile$1$ [26]),
    .i10(\t/a/regfile/regfile$10$ [26]),
    .i11(\t/a/regfile/regfile$11$ [26]),
    .i12(\t/a/regfile/regfile$12$ [26]),
    .i13(\t/a/regfile/regfile$13$ [26]),
    .i14(\t/a/regfile/regfile$14$ [26]),
    .i15(\t/a/regfile/regfile$15$ [26]),
    .i16(\t/a/regfile/regfile$16$ [26]),
    .i17(\t/a/regfile/regfile$17$ [26]),
    .i18(\t/a/regfile/regfile$18$ [26]),
    .i19(\t/a/regfile/regfile$19$ [26]),
    .i2(\t/a/regfile/regfile$2$ [26]),
    .i20(\t/a/regfile/regfile$20$ [26]),
    .i21(\t/a/regfile/regfile$21$ [26]),
    .i22(\t/a/regfile/regfile$22$ [26]),
    .i23(\t/a/regfile/regfile$23$ [26]),
    .i24(\t/a/regfile/regfile$24$ [26]),
    .i25(\t/a/regfile/regfile$25$ [26]),
    .i26(\t/a/regfile/regfile$26$ [26]),
    .i27(\t/a/regfile/regfile$27$ [26]),
    .i28(\t/a/regfile/regfile$28$ [26]),
    .i29(\t/a/regfile/regfile$29$ [26]),
    .i3(\t/a/regfile/regfile$3$ [26]),
    .i30(\t/a/regfile/regfile$30$ [26]),
    .i31(\t/a/regfile/regfile$31$ [26]),
    .i4(\t/a/regfile/regfile$4$ [26]),
    .i5(\t/a/regfile/regfile$5$ [26]),
    .i6(\t/a/regfile/regfile$6$ [26]),
    .i7(\t/a/regfile/regfile$7$ [26]),
    .i8(\t/a/regfile/regfile$8$ [26]),
    .i9(\t/a/regfile/regfile$9$ [26]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [26]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b27  (
    .i0(\t/a/regfile/regfile$0$ [27]),
    .i1(\t/a/regfile/regfile$1$ [27]),
    .i10(\t/a/regfile/regfile$10$ [27]),
    .i11(\t/a/regfile/regfile$11$ [27]),
    .i12(\t/a/regfile/regfile$12$ [27]),
    .i13(\t/a/regfile/regfile$13$ [27]),
    .i14(\t/a/regfile/regfile$14$ [27]),
    .i15(\t/a/regfile/regfile$15$ [27]),
    .i16(\t/a/regfile/regfile$16$ [27]),
    .i17(\t/a/regfile/regfile$17$ [27]),
    .i18(\t/a/regfile/regfile$18$ [27]),
    .i19(\t/a/regfile/regfile$19$ [27]),
    .i2(\t/a/regfile/regfile$2$ [27]),
    .i20(\t/a/regfile/regfile$20$ [27]),
    .i21(\t/a/regfile/regfile$21$ [27]),
    .i22(\t/a/regfile/regfile$22$ [27]),
    .i23(\t/a/regfile/regfile$23$ [27]),
    .i24(\t/a/regfile/regfile$24$ [27]),
    .i25(\t/a/regfile/regfile$25$ [27]),
    .i26(\t/a/regfile/regfile$26$ [27]),
    .i27(\t/a/regfile/regfile$27$ [27]),
    .i28(\t/a/regfile/regfile$28$ [27]),
    .i29(\t/a/regfile/regfile$29$ [27]),
    .i3(\t/a/regfile/regfile$3$ [27]),
    .i30(\t/a/regfile/regfile$30$ [27]),
    .i31(\t/a/regfile/regfile$31$ [27]),
    .i4(\t/a/regfile/regfile$4$ [27]),
    .i5(\t/a/regfile/regfile$5$ [27]),
    .i6(\t/a/regfile/regfile$6$ [27]),
    .i7(\t/a/regfile/regfile$7$ [27]),
    .i8(\t/a/regfile/regfile$8$ [27]),
    .i9(\t/a/regfile/regfile$9$ [27]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [27]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b28  (
    .i0(\t/a/regfile/regfile$0$ [28]),
    .i1(\t/a/regfile/regfile$1$ [28]),
    .i10(\t/a/regfile/regfile$10$ [28]),
    .i11(\t/a/regfile/regfile$11$ [28]),
    .i12(\t/a/regfile/regfile$12$ [28]),
    .i13(\t/a/regfile/regfile$13$ [28]),
    .i14(\t/a/regfile/regfile$14$ [28]),
    .i15(\t/a/regfile/regfile$15$ [28]),
    .i16(\t/a/regfile/regfile$16$ [28]),
    .i17(\t/a/regfile/regfile$17$ [28]),
    .i18(\t/a/regfile/regfile$18$ [28]),
    .i19(\t/a/regfile/regfile$19$ [28]),
    .i2(\t/a/regfile/regfile$2$ [28]),
    .i20(\t/a/regfile/regfile$20$ [28]),
    .i21(\t/a/regfile/regfile$21$ [28]),
    .i22(\t/a/regfile/regfile$22$ [28]),
    .i23(\t/a/regfile/regfile$23$ [28]),
    .i24(\t/a/regfile/regfile$24$ [28]),
    .i25(\t/a/regfile/regfile$25$ [28]),
    .i26(\t/a/regfile/regfile$26$ [28]),
    .i27(\t/a/regfile/regfile$27$ [28]),
    .i28(\t/a/regfile/regfile$28$ [28]),
    .i29(\t/a/regfile/regfile$29$ [28]),
    .i3(\t/a/regfile/regfile$3$ [28]),
    .i30(\t/a/regfile/regfile$30$ [28]),
    .i31(\t/a/regfile/regfile$31$ [28]),
    .i4(\t/a/regfile/regfile$4$ [28]),
    .i5(\t/a/regfile/regfile$5$ [28]),
    .i6(\t/a/regfile/regfile$6$ [28]),
    .i7(\t/a/regfile/regfile$7$ [28]),
    .i8(\t/a/regfile/regfile$8$ [28]),
    .i9(\t/a/regfile/regfile$9$ [28]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [28]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b29  (
    .i0(\t/a/regfile/regfile$0$ [29]),
    .i1(\t/a/regfile/regfile$1$ [29]),
    .i10(\t/a/regfile/regfile$10$ [29]),
    .i11(\t/a/regfile/regfile$11$ [29]),
    .i12(\t/a/regfile/regfile$12$ [29]),
    .i13(\t/a/regfile/regfile$13$ [29]),
    .i14(\t/a/regfile/regfile$14$ [29]),
    .i15(\t/a/regfile/regfile$15$ [29]),
    .i16(\t/a/regfile/regfile$16$ [29]),
    .i17(\t/a/regfile/regfile$17$ [29]),
    .i18(\t/a/regfile/regfile$18$ [29]),
    .i19(\t/a/regfile/regfile$19$ [29]),
    .i2(\t/a/regfile/regfile$2$ [29]),
    .i20(\t/a/regfile/regfile$20$ [29]),
    .i21(\t/a/regfile/regfile$21$ [29]),
    .i22(\t/a/regfile/regfile$22$ [29]),
    .i23(\t/a/regfile/regfile$23$ [29]),
    .i24(\t/a/regfile/regfile$24$ [29]),
    .i25(\t/a/regfile/regfile$25$ [29]),
    .i26(\t/a/regfile/regfile$26$ [29]),
    .i27(\t/a/regfile/regfile$27$ [29]),
    .i28(\t/a/regfile/regfile$28$ [29]),
    .i29(\t/a/regfile/regfile$29$ [29]),
    .i3(\t/a/regfile/regfile$3$ [29]),
    .i30(\t/a/regfile/regfile$30$ [29]),
    .i31(\t/a/regfile/regfile$31$ [29]),
    .i4(\t/a/regfile/regfile$4$ [29]),
    .i5(\t/a/regfile/regfile$5$ [29]),
    .i6(\t/a/regfile/regfile$6$ [29]),
    .i7(\t/a/regfile/regfile$7$ [29]),
    .i8(\t/a/regfile/regfile$8$ [29]),
    .i9(\t/a/regfile/regfile$9$ [29]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [29]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b3  (
    .i0(\t/a/regfile/regfile$0$ [3]),
    .i1(\t/a/regfile/regfile$1$ [3]),
    .i10(\t/a/regfile/regfile$10$ [3]),
    .i11(\t/a/regfile/regfile$11$ [3]),
    .i12(\t/a/regfile/regfile$12$ [3]),
    .i13(\t/a/regfile/regfile$13$ [3]),
    .i14(\t/a/regfile/regfile$14$ [3]),
    .i15(\t/a/regfile/regfile$15$ [3]),
    .i16(\t/a/regfile/regfile$16$ [3]),
    .i17(\t/a/regfile/regfile$17$ [3]),
    .i18(\t/a/regfile/regfile$18$ [3]),
    .i19(\t/a/regfile/regfile$19$ [3]),
    .i2(\t/a/regfile/regfile$2$ [3]),
    .i20(\t/a/regfile/regfile$20$ [3]),
    .i21(\t/a/regfile/regfile$21$ [3]),
    .i22(\t/a/regfile/regfile$22$ [3]),
    .i23(\t/a/regfile/regfile$23$ [3]),
    .i24(\t/a/regfile/regfile$24$ [3]),
    .i25(\t/a/regfile/regfile$25$ [3]),
    .i26(\t/a/regfile/regfile$26$ [3]),
    .i27(\t/a/regfile/regfile$27$ [3]),
    .i28(\t/a/regfile/regfile$28$ [3]),
    .i29(\t/a/regfile/regfile$29$ [3]),
    .i3(\t/a/regfile/regfile$3$ [3]),
    .i30(\t/a/regfile/regfile$30$ [3]),
    .i31(\t/a/regfile/regfile$31$ [3]),
    .i4(\t/a/regfile/regfile$4$ [3]),
    .i5(\t/a/regfile/regfile$5$ [3]),
    .i6(\t/a/regfile/regfile$6$ [3]),
    .i7(\t/a/regfile/regfile$7$ [3]),
    .i8(\t/a/regfile/regfile$8$ [3]),
    .i9(\t/a/regfile/regfile$9$ [3]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [3]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b30  (
    .i0(\t/a/regfile/regfile$0$ [30]),
    .i1(\t/a/regfile/regfile$1$ [30]),
    .i10(\t/a/regfile/regfile$10$ [30]),
    .i11(\t/a/regfile/regfile$11$ [30]),
    .i12(\t/a/regfile/regfile$12$ [30]),
    .i13(\t/a/regfile/regfile$13$ [30]),
    .i14(\t/a/regfile/regfile$14$ [30]),
    .i15(\t/a/regfile/regfile$15$ [30]),
    .i16(\t/a/regfile/regfile$16$ [30]),
    .i17(\t/a/regfile/regfile$17$ [30]),
    .i18(\t/a/regfile/regfile$18$ [30]),
    .i19(\t/a/regfile/regfile$19$ [30]),
    .i2(\t/a/regfile/regfile$2$ [30]),
    .i20(\t/a/regfile/regfile$20$ [30]),
    .i21(\t/a/regfile/regfile$21$ [30]),
    .i22(\t/a/regfile/regfile$22$ [30]),
    .i23(\t/a/regfile/regfile$23$ [30]),
    .i24(\t/a/regfile/regfile$24$ [30]),
    .i25(\t/a/regfile/regfile$25$ [30]),
    .i26(\t/a/regfile/regfile$26$ [30]),
    .i27(\t/a/regfile/regfile$27$ [30]),
    .i28(\t/a/regfile/regfile$28$ [30]),
    .i29(\t/a/regfile/regfile$29$ [30]),
    .i3(\t/a/regfile/regfile$3$ [30]),
    .i30(\t/a/regfile/regfile$30$ [30]),
    .i31(\t/a/regfile/regfile$31$ [30]),
    .i4(\t/a/regfile/regfile$4$ [30]),
    .i5(\t/a/regfile/regfile$5$ [30]),
    .i6(\t/a/regfile/regfile$6$ [30]),
    .i7(\t/a/regfile/regfile$7$ [30]),
    .i8(\t/a/regfile/regfile$8$ [30]),
    .i9(\t/a/regfile/regfile$9$ [30]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [30]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b31  (
    .i0(\t/a/regfile/regfile$0$ [31]),
    .i1(\t/a/regfile/regfile$1$ [31]),
    .i10(\t/a/regfile/regfile$10$ [31]),
    .i11(\t/a/regfile/regfile$11$ [31]),
    .i12(\t/a/regfile/regfile$12$ [31]),
    .i13(\t/a/regfile/regfile$13$ [31]),
    .i14(\t/a/regfile/regfile$14$ [31]),
    .i15(\t/a/regfile/regfile$15$ [31]),
    .i16(\t/a/regfile/regfile$16$ [31]),
    .i17(\t/a/regfile/regfile$17$ [31]),
    .i18(\t/a/regfile/regfile$18$ [31]),
    .i19(\t/a/regfile/regfile$19$ [31]),
    .i2(\t/a/regfile/regfile$2$ [31]),
    .i20(\t/a/regfile/regfile$20$ [31]),
    .i21(\t/a/regfile/regfile$21$ [31]),
    .i22(\t/a/regfile/regfile$22$ [31]),
    .i23(\t/a/regfile/regfile$23$ [31]),
    .i24(\t/a/regfile/regfile$24$ [31]),
    .i25(\t/a/regfile/regfile$25$ [31]),
    .i26(\t/a/regfile/regfile$26$ [31]),
    .i27(\t/a/regfile/regfile$27$ [31]),
    .i28(\t/a/regfile/regfile$28$ [31]),
    .i29(\t/a/regfile/regfile$29$ [31]),
    .i3(\t/a/regfile/regfile$3$ [31]),
    .i30(\t/a/regfile/regfile$30$ [31]),
    .i31(\t/a/regfile/regfile$31$ [31]),
    .i4(\t/a/regfile/regfile$4$ [31]),
    .i5(\t/a/regfile/regfile$5$ [31]),
    .i6(\t/a/regfile/regfile$6$ [31]),
    .i7(\t/a/regfile/regfile$7$ [31]),
    .i8(\t/a/regfile/regfile$8$ [31]),
    .i9(\t/a/regfile/regfile$9$ [31]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n7 [31]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b36  (
    .i0(\t/a/regfile/regfile$0$ [4]),
    .i1(\t/a/regfile/regfile$1$ [4]),
    .i10(\t/a/regfile/regfile$10$ [4]),
    .i11(\t/a/regfile/regfile$11$ [4]),
    .i12(\t/a/regfile/regfile$12$ [4]),
    .i13(\t/a/regfile/regfile$13$ [4]),
    .i14(\t/a/regfile/regfile$14$ [4]),
    .i15(\t/a/regfile/regfile$15$ [4]),
    .i16(\t/a/regfile/regfile$16$ [4]),
    .i17(\t/a/regfile/regfile$17$ [4]),
    .i18(\t/a/regfile/regfile$18$ [4]),
    .i19(\t/a/regfile/regfile$19$ [4]),
    .i2(\t/a/regfile/regfile$2$ [4]),
    .i20(\t/a/regfile/regfile$20$ [4]),
    .i21(\t/a/regfile/regfile$21$ [4]),
    .i22(\t/a/regfile/regfile$22$ [4]),
    .i23(\t/a/regfile/regfile$23$ [4]),
    .i24(\t/a/regfile/regfile$24$ [4]),
    .i25(\t/a/regfile/regfile$25$ [4]),
    .i26(\t/a/regfile/regfile$26$ [4]),
    .i27(\t/a/regfile/regfile$27$ [4]),
    .i28(\t/a/regfile/regfile$28$ [4]),
    .i29(\t/a/regfile/regfile$29$ [4]),
    .i3(\t/a/regfile/regfile$3$ [4]),
    .i30(\t/a/regfile/regfile$30$ [4]),
    .i31(\t/a/regfile/regfile$31$ [4]),
    .i4(\t/a/regfile/regfile$4$ [4]),
    .i5(\t/a/regfile/regfile$5$ [4]),
    .i6(\t/a/regfile/regfile$6$ [4]),
    .i7(\t/a/regfile/regfile$7$ [4]),
    .i8(\t/a/regfile/regfile$8$ [4]),
    .i9(\t/a/regfile/regfile$9$ [4]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n8 [4]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b37  (
    .i0(\t/a/regfile/regfile$0$ [5]),
    .i1(\t/a/regfile/regfile$1$ [5]),
    .i10(\t/a/regfile/regfile$10$ [5]),
    .i11(\t/a/regfile/regfile$11$ [5]),
    .i12(\t/a/regfile/regfile$12$ [5]),
    .i13(\t/a/regfile/regfile$13$ [5]),
    .i14(\t/a/regfile/regfile$14$ [5]),
    .i15(\t/a/regfile/regfile$15$ [5]),
    .i16(\t/a/regfile/regfile$16$ [5]),
    .i17(\t/a/regfile/regfile$17$ [5]),
    .i18(\t/a/regfile/regfile$18$ [5]),
    .i19(\t/a/regfile/regfile$19$ [5]),
    .i2(\t/a/regfile/regfile$2$ [5]),
    .i20(\t/a/regfile/regfile$20$ [5]),
    .i21(\t/a/regfile/regfile$21$ [5]),
    .i22(\t/a/regfile/regfile$22$ [5]),
    .i23(\t/a/regfile/regfile$23$ [5]),
    .i24(\t/a/regfile/regfile$24$ [5]),
    .i25(\t/a/regfile/regfile$25$ [5]),
    .i26(\t/a/regfile/regfile$26$ [5]),
    .i27(\t/a/regfile/regfile$27$ [5]),
    .i28(\t/a/regfile/regfile$28$ [5]),
    .i29(\t/a/regfile/regfile$29$ [5]),
    .i3(\t/a/regfile/regfile$3$ [5]),
    .i30(\t/a/regfile/regfile$30$ [5]),
    .i31(\t/a/regfile/regfile$31$ [5]),
    .i4(\t/a/regfile/regfile$4$ [5]),
    .i5(\t/a/regfile/regfile$5$ [5]),
    .i6(\t/a/regfile/regfile$6$ [5]),
    .i7(\t/a/regfile/regfile$7$ [5]),
    .i8(\t/a/regfile/regfile$8$ [5]),
    .i9(\t/a/regfile/regfile$9$ [5]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n8 [5]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b38  (
    .i0(\t/a/regfile/regfile$0$ [6]),
    .i1(\t/a/regfile/regfile$1$ [6]),
    .i10(\t/a/regfile/regfile$10$ [6]),
    .i11(\t/a/regfile/regfile$11$ [6]),
    .i12(\t/a/regfile/regfile$12$ [6]),
    .i13(\t/a/regfile/regfile$13$ [6]),
    .i14(\t/a/regfile/regfile$14$ [6]),
    .i15(\t/a/regfile/regfile$15$ [6]),
    .i16(\t/a/regfile/regfile$16$ [6]),
    .i17(\t/a/regfile/regfile$17$ [6]),
    .i18(\t/a/regfile/regfile$18$ [6]),
    .i19(\t/a/regfile/regfile$19$ [6]),
    .i2(\t/a/regfile/regfile$2$ [6]),
    .i20(\t/a/regfile/regfile$20$ [6]),
    .i21(\t/a/regfile/regfile$21$ [6]),
    .i22(\t/a/regfile/regfile$22$ [6]),
    .i23(\t/a/regfile/regfile$23$ [6]),
    .i24(\t/a/regfile/regfile$24$ [6]),
    .i25(\t/a/regfile/regfile$25$ [6]),
    .i26(\t/a/regfile/regfile$26$ [6]),
    .i27(\t/a/regfile/regfile$27$ [6]),
    .i28(\t/a/regfile/regfile$28$ [6]),
    .i29(\t/a/regfile/regfile$29$ [6]),
    .i3(\t/a/regfile/regfile$3$ [6]),
    .i30(\t/a/regfile/regfile$30$ [6]),
    .i31(\t/a/regfile/regfile$31$ [6]),
    .i4(\t/a/regfile/regfile$4$ [6]),
    .i5(\t/a/regfile/regfile$5$ [6]),
    .i6(\t/a/regfile/regfile$6$ [6]),
    .i7(\t/a/regfile/regfile$7$ [6]),
    .i8(\t/a/regfile/regfile$8$ [6]),
    .i9(\t/a/regfile/regfile$9$ [6]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n8 [6]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b39  (
    .i0(\t/a/regfile/regfile$0$ [7]),
    .i1(\t/a/regfile/regfile$1$ [7]),
    .i10(\t/a/regfile/regfile$10$ [7]),
    .i11(\t/a/regfile/regfile$11$ [7]),
    .i12(\t/a/regfile/regfile$12$ [7]),
    .i13(\t/a/regfile/regfile$13$ [7]),
    .i14(\t/a/regfile/regfile$14$ [7]),
    .i15(\t/a/regfile/regfile$15$ [7]),
    .i16(\t/a/regfile/regfile$16$ [7]),
    .i17(\t/a/regfile/regfile$17$ [7]),
    .i18(\t/a/regfile/regfile$18$ [7]),
    .i19(\t/a/regfile/regfile$19$ [7]),
    .i2(\t/a/regfile/regfile$2$ [7]),
    .i20(\t/a/regfile/regfile$20$ [7]),
    .i21(\t/a/regfile/regfile$21$ [7]),
    .i22(\t/a/regfile/regfile$22$ [7]),
    .i23(\t/a/regfile/regfile$23$ [7]),
    .i24(\t/a/regfile/regfile$24$ [7]),
    .i25(\t/a/regfile/regfile$25$ [7]),
    .i26(\t/a/regfile/regfile$26$ [7]),
    .i27(\t/a/regfile/regfile$27$ [7]),
    .i28(\t/a/regfile/regfile$28$ [7]),
    .i29(\t/a/regfile/regfile$29$ [7]),
    .i3(\t/a/regfile/regfile$3$ [7]),
    .i30(\t/a/regfile/regfile$30$ [7]),
    .i31(\t/a/regfile/regfile$31$ [7]),
    .i4(\t/a/regfile/regfile$4$ [7]),
    .i5(\t/a/regfile/regfile$5$ [7]),
    .i6(\t/a/regfile/regfile$6$ [7]),
    .i7(\t/a/regfile/regfile$7$ [7]),
    .i8(\t/a/regfile/regfile$8$ [7]),
    .i9(\t/a/regfile/regfile$9$ [7]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n8 [7]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b40  (
    .i0(\t/a/regfile/regfile$0$ [8]),
    .i1(\t/a/regfile/regfile$1$ [8]),
    .i10(\t/a/regfile/regfile$10$ [8]),
    .i11(\t/a/regfile/regfile$11$ [8]),
    .i12(\t/a/regfile/regfile$12$ [8]),
    .i13(\t/a/regfile/regfile$13$ [8]),
    .i14(\t/a/regfile/regfile$14$ [8]),
    .i15(\t/a/regfile/regfile$15$ [8]),
    .i16(\t/a/regfile/regfile$16$ [8]),
    .i17(\t/a/regfile/regfile$17$ [8]),
    .i18(\t/a/regfile/regfile$18$ [8]),
    .i19(\t/a/regfile/regfile$19$ [8]),
    .i2(\t/a/regfile/regfile$2$ [8]),
    .i20(\t/a/regfile/regfile$20$ [8]),
    .i21(\t/a/regfile/regfile$21$ [8]),
    .i22(\t/a/regfile/regfile$22$ [8]),
    .i23(\t/a/regfile/regfile$23$ [8]),
    .i24(\t/a/regfile/regfile$24$ [8]),
    .i25(\t/a/regfile/regfile$25$ [8]),
    .i26(\t/a/regfile/regfile$26$ [8]),
    .i27(\t/a/regfile/regfile$27$ [8]),
    .i28(\t/a/regfile/regfile$28$ [8]),
    .i29(\t/a/regfile/regfile$29$ [8]),
    .i3(\t/a/regfile/regfile$3$ [8]),
    .i30(\t/a/regfile/regfile$30$ [8]),
    .i31(\t/a/regfile/regfile$31$ [8]),
    .i4(\t/a/regfile/regfile$4$ [8]),
    .i5(\t/a/regfile/regfile$5$ [8]),
    .i6(\t/a/regfile/regfile$6$ [8]),
    .i7(\t/a/regfile/regfile$7$ [8]),
    .i8(\t/a/regfile/regfile$8$ [8]),
    .i9(\t/a/regfile/regfile$9$ [8]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n8 [8]));  // register.v(23)
  binary_mux_s5_w1 \t/a/regfile/mux40_b41  (
    .i0(\t/a/regfile/regfile$0$ [9]),
    .i1(\t/a/regfile/regfile$1$ [9]),
    .i10(\t/a/regfile/regfile$10$ [9]),
    .i11(\t/a/regfile/regfile$11$ [9]),
    .i12(\t/a/regfile/regfile$12$ [9]),
    .i13(\t/a/regfile/regfile$13$ [9]),
    .i14(\t/a/regfile/regfile$14$ [9]),
    .i15(\t/a/regfile/regfile$15$ [9]),
    .i16(\t/a/regfile/regfile$16$ [9]),
    .i17(\t/a/regfile/regfile$17$ [9]),
    .i18(\t/a/regfile/regfile$18$ [9]),
    .i19(\t/a/regfile/regfile$19$ [9]),
    .i2(\t/a/regfile/regfile$2$ [9]),
    .i20(\t/a/regfile/regfile$20$ [9]),
    .i21(\t/a/regfile/regfile$21$ [9]),
    .i22(\t/a/regfile/regfile$22$ [9]),
    .i23(\t/a/regfile/regfile$23$ [9]),
    .i24(\t/a/regfile/regfile$24$ [9]),
    .i25(\t/a/regfile/regfile$25$ [9]),
    .i26(\t/a/regfile/regfile$26$ [9]),
    .i27(\t/a/regfile/regfile$27$ [9]),
    .i28(\t/a/regfile/regfile$28$ [9]),
    .i29(\t/a/regfile/regfile$29$ [9]),
    .i3(\t/a/regfile/regfile$3$ [9]),
    .i30(\t/a/regfile/regfile$30$ [9]),
    .i31(\t/a/regfile/regfile$31$ [9]),
    .i4(\t/a/regfile/regfile$4$ [9]),
    .i5(\t/a/regfile/regfile$5$ [9]),
    .i6(\t/a/regfile/regfile$6$ [9]),
    .i7(\t/a/regfile/regfile$7$ [9]),
    .i8(\t/a/regfile/regfile$8$ [9]),
    .i9(\t/a/regfile/regfile$9$ [9]),
    .sel(\t/a/ID_rs1 ),
    .o(\t/a/regfile/n8 [9]));  // register.v(23)
  and \t/a/regfile/mux4_b0_sel_is_2  (\t/a/regfile/mux4_b0_sel_is_2_o , \t/a/regfile/n2_neg , \t/a/regfile/n6 );
  not \t/a/regfile/mux4_b0_sel_is_2_o_inv  (\t/a/regfile/mux4_b0_sel_is_2_o_neg , \t/a/regfile/mux4_b0_sel_is_2_o );
  AL_MUX \t/a/regfile/mux5_b0  (
    .i0(\t/a/reg_writedat [0]),
    .i1(\t/a/regfile/n7 [0]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [0]));
  and \t/a/regfile/mux5_b0_sel_is_0  (\t/a/regfile/mux5_b0_sel_is_0_o , \t/a/regfile/n4_neg , \t/a/regfile/n2_neg );
  AL_MUX \t/a/regfile/mux5_b1  (
    .i0(\t/a/reg_writedat [1]),
    .i1(\t/a/regfile/n7 [1]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [1]));
  AL_MUX \t/a/regfile/mux5_b10  (
    .i0(\t/a/reg_writedat [10]),
    .i1(\t/a/regfile/n7 [10]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [10]));
  AL_MUX \t/a/regfile/mux5_b11  (
    .i0(\t/a/reg_writedat [11]),
    .i1(\t/a/regfile/n7 [11]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [11]));
  AL_MUX \t/a/regfile/mux5_b12  (
    .i0(\t/a/reg_writedat [12]),
    .i1(\t/a/regfile/n7 [12]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [12]));
  AL_MUX \t/a/regfile/mux5_b13  (
    .i0(\t/a/reg_writedat [13]),
    .i1(\t/a/regfile/n7 [13]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [13]));
  AL_MUX \t/a/regfile/mux5_b14  (
    .i0(\t/a/reg_writedat [14]),
    .i1(\t/a/regfile/n7 [14]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [14]));
  AL_MUX \t/a/regfile/mux5_b15  (
    .i0(\t/a/reg_writedat [15]),
    .i1(\t/a/regfile/n7 [15]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [15]));
  AL_MUX \t/a/regfile/mux5_b16  (
    .i0(\t/a/reg_writedat [16]),
    .i1(\t/a/regfile/n7 [16]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [16]));
  AL_MUX \t/a/regfile/mux5_b17  (
    .i0(\t/a/reg_writedat [17]),
    .i1(\t/a/regfile/n7 [17]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [17]));
  AL_MUX \t/a/regfile/mux5_b18  (
    .i0(\t/a/reg_writedat [18]),
    .i1(\t/a/regfile/n7 [18]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [18]));
  AL_MUX \t/a/regfile/mux5_b19  (
    .i0(\t/a/reg_writedat [19]),
    .i1(\t/a/regfile/n7 [19]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [19]));
  AL_MUX \t/a/regfile/mux5_b2  (
    .i0(\t/a/reg_writedat [2]),
    .i1(\t/a/regfile/n7 [2]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [2]));
  AL_MUX \t/a/regfile/mux5_b20  (
    .i0(\t/a/reg_writedat [20]),
    .i1(\t/a/regfile/n7 [20]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [20]));
  AL_MUX \t/a/regfile/mux5_b21  (
    .i0(\t/a/reg_writedat [21]),
    .i1(\t/a/regfile/n7 [21]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [21]));
  AL_MUX \t/a/regfile/mux5_b22  (
    .i0(\t/a/reg_writedat [22]),
    .i1(\t/a/regfile/n7 [22]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [22]));
  AL_MUX \t/a/regfile/mux5_b23  (
    .i0(\t/a/reg_writedat [23]),
    .i1(\t/a/regfile/n7 [23]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [23]));
  AL_MUX \t/a/regfile/mux5_b24  (
    .i0(\t/a/reg_writedat [24]),
    .i1(\t/a/regfile/n7 [24]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [24]));
  AL_MUX \t/a/regfile/mux5_b25  (
    .i0(\t/a/reg_writedat [25]),
    .i1(\t/a/regfile/n7 [25]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [25]));
  AL_MUX \t/a/regfile/mux5_b26  (
    .i0(\t/a/reg_writedat [26]),
    .i1(\t/a/regfile/n7 [26]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [26]));
  AL_MUX \t/a/regfile/mux5_b27  (
    .i0(\t/a/reg_writedat [27]),
    .i1(\t/a/regfile/n7 [27]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [27]));
  AL_MUX \t/a/regfile/mux5_b28  (
    .i0(\t/a/reg_writedat [28]),
    .i1(\t/a/regfile/n7 [28]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [28]));
  AL_MUX \t/a/regfile/mux5_b29  (
    .i0(\t/a/reg_writedat [29]),
    .i1(\t/a/regfile/n7 [29]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [29]));
  AL_MUX \t/a/regfile/mux5_b3  (
    .i0(\t/a/reg_writedat [3]),
    .i1(\t/a/regfile/n7 [3]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [3]));
  AL_MUX \t/a/regfile/mux5_b30  (
    .i0(\t/a/reg_writedat [30]),
    .i1(\t/a/regfile/n7 [30]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [30]));
  AL_MUX \t/a/regfile/mux5_b31  (
    .i0(\t/a/reg_writedat [31]),
    .i1(\t/a/regfile/n7 [31]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [31]));
  AL_MUX \t/a/regfile/mux5_b4  (
    .i0(\t/a/reg_writedat [4]),
    .i1(\t/a/regfile/n8 [4]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [4]));
  AL_MUX \t/a/regfile/mux5_b5  (
    .i0(\t/a/reg_writedat [5]),
    .i1(\t/a/regfile/n8 [5]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [5]));
  AL_MUX \t/a/regfile/mux5_b6  (
    .i0(\t/a/reg_writedat [6]),
    .i1(\t/a/regfile/n8 [6]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [6]));
  AL_MUX \t/a/regfile/mux5_b7  (
    .i0(\t/a/reg_writedat [7]),
    .i1(\t/a/regfile/n8 [7]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [7]));
  AL_MUX \t/a/regfile/mux5_b8  (
    .i0(\t/a/reg_writedat [8]),
    .i1(\t/a/regfile/n8 [8]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [8]));
  AL_MUX \t/a/regfile/mux5_b9  (
    .i0(\t/a/reg_writedat [9]),
    .i1(\t/a/regfile/n8 [9]),
    .sel(\t/a/regfile/mux5_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat1 [9]));
  AL_MUX \t/a/regfile/mux6_b0  (
    .i0(\t/a/reg_writedat [0]),
    .i1(\t/a/regfile/n5 [0]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [0]));
  and \t/a/regfile/mux6_b0_sel_is_0  (\t/a/regfile/mux6_b0_sel_is_0_o , \t/a/regfile/n4_neg , \t/a/regfile/mux4_b0_sel_is_2_o_neg );
  AL_MUX \t/a/regfile/mux6_b1  (
    .i0(\t/a/reg_writedat [1]),
    .i1(\t/a/regfile/n5 [1]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [1]));
  AL_MUX \t/a/regfile/mux6_b10  (
    .i0(\t/a/reg_writedat [10]),
    .i1(\t/a/regfile/n5 [10]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [10]));
  AL_MUX \t/a/regfile/mux6_b11  (
    .i0(\t/a/reg_writedat [11]),
    .i1(\t/a/regfile/n5 [11]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [11]));
  AL_MUX \t/a/regfile/mux6_b12  (
    .i0(\t/a/reg_writedat [12]),
    .i1(\t/a/regfile/n5 [12]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [12]));
  AL_MUX \t/a/regfile/mux6_b13  (
    .i0(\t/a/reg_writedat [13]),
    .i1(\t/a/regfile/n5 [13]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [13]));
  AL_MUX \t/a/regfile/mux6_b14  (
    .i0(\t/a/reg_writedat [14]),
    .i1(\t/a/regfile/n5 [14]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [14]));
  AL_MUX \t/a/regfile/mux6_b15  (
    .i0(\t/a/reg_writedat [15]),
    .i1(\t/a/regfile/n5 [15]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [15]));
  AL_MUX \t/a/regfile/mux6_b16  (
    .i0(\t/a/reg_writedat [16]),
    .i1(\t/a/regfile/n5 [16]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [16]));
  AL_MUX \t/a/regfile/mux6_b17  (
    .i0(\t/a/reg_writedat [17]),
    .i1(\t/a/regfile/n5 [17]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [17]));
  AL_MUX \t/a/regfile/mux6_b18  (
    .i0(\t/a/reg_writedat [18]),
    .i1(\t/a/regfile/n5 [18]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [18]));
  AL_MUX \t/a/regfile/mux6_b19  (
    .i0(\t/a/reg_writedat [19]),
    .i1(\t/a/regfile/n5 [19]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [19]));
  AL_MUX \t/a/regfile/mux6_b2  (
    .i0(\t/a/reg_writedat [2]),
    .i1(\t/a/regfile/n5 [2]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [2]));
  AL_MUX \t/a/regfile/mux6_b20  (
    .i0(\t/a/reg_writedat [20]),
    .i1(\t/a/regfile/n5 [20]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [20]));
  AL_MUX \t/a/regfile/mux6_b21  (
    .i0(\t/a/reg_writedat [21]),
    .i1(\t/a/regfile/n5 [21]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [21]));
  AL_MUX \t/a/regfile/mux6_b22  (
    .i0(\t/a/reg_writedat [22]),
    .i1(\t/a/regfile/n5 [22]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [22]));
  AL_MUX \t/a/regfile/mux6_b23  (
    .i0(\t/a/reg_writedat [23]),
    .i1(\t/a/regfile/n5 [23]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [23]));
  AL_MUX \t/a/regfile/mux6_b24  (
    .i0(\t/a/reg_writedat [24]),
    .i1(\t/a/regfile/n5 [24]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [24]));
  AL_MUX \t/a/regfile/mux6_b25  (
    .i0(\t/a/reg_writedat [25]),
    .i1(\t/a/regfile/n5 [25]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [25]));
  AL_MUX \t/a/regfile/mux6_b26  (
    .i0(\t/a/reg_writedat [26]),
    .i1(\t/a/regfile/n5 [26]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [26]));
  AL_MUX \t/a/regfile/mux6_b27  (
    .i0(\t/a/reg_writedat [27]),
    .i1(\t/a/regfile/n5 [27]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [27]));
  AL_MUX \t/a/regfile/mux6_b28  (
    .i0(\t/a/reg_writedat [28]),
    .i1(\t/a/regfile/n5 [28]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [28]));
  AL_MUX \t/a/regfile/mux6_b29  (
    .i0(\t/a/reg_writedat [29]),
    .i1(\t/a/regfile/n5 [29]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [29]));
  AL_MUX \t/a/regfile/mux6_b3  (
    .i0(\t/a/reg_writedat [3]),
    .i1(\t/a/regfile/n5 [3]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [3]));
  AL_MUX \t/a/regfile/mux6_b30  (
    .i0(\t/a/reg_writedat [30]),
    .i1(\t/a/regfile/n5 [30]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [30]));
  AL_MUX \t/a/regfile/mux6_b31  (
    .i0(\t/a/reg_writedat [31]),
    .i1(\t/a/regfile/n5 [31]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [31]));
  AL_MUX \t/a/regfile/mux6_b4  (
    .i0(\t/a/reg_writedat [4]),
    .i1(\t/a/regfile/n5 [4]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [4]));
  AL_MUX \t/a/regfile/mux6_b5  (
    .i0(\t/a/reg_writedat [5]),
    .i1(\t/a/regfile/n5 [5]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [5]));
  AL_MUX \t/a/regfile/mux6_b6  (
    .i0(\t/a/reg_writedat [6]),
    .i1(\t/a/regfile/n5 [6]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [6]));
  AL_MUX \t/a/regfile/mux6_b7  (
    .i0(\t/a/reg_writedat [7]),
    .i1(\t/a/regfile/n5 [7]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [7]));
  AL_MUX \t/a/regfile/mux6_b8  (
    .i0(\t/a/reg_writedat [8]),
    .i1(\t/a/regfile/n5 [8]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [8]));
  AL_MUX \t/a/regfile/mux6_b9  (
    .i0(\t/a/reg_writedat [9]),
    .i1(\t/a/regfile/n5 [9]),
    .sel(\t/a/regfile/mux6_b0_sel_is_0_o ),
    .o(\t/a/ID_read_dat2 [9]));
  not \t/a/regfile/n2_inv  (\t/a/regfile/n2_neg , \t/a/regfile/n2 );
  not \t/a/regfile/n4_inv  (\t/a/regfile/n4_neg , \t/a/regfile/n4 );
  reg_ar_as_w1 \t/a/regfile/reg0_b0  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b10  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b100  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1000  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1001  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1002  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1003  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1004  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1005  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1006  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1007  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1008  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1009  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b101  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$3$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1010  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1011  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1012  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1013  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1014  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1015  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1016  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1017  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1018  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1019  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b102  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1020  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1021  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1022  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b1023  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b103  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b104  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b105  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b106  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b107  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b108  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b109  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b11  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b110  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b111  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b112  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b113  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b114  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b115  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b116  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b117  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b118  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b119  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b12  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b120  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b121  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b122  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b123  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b124  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b125  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b126  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b127  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b128  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$4$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b129  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b13  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b130  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$4$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b131  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b132  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$4$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b133  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b134  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b135  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b136  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b137  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b138  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b139  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b14  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b140  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b141  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b142  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b143  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b144  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b145  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b146  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b147  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b148  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b149  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b15  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b150  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b151  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b152  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b153  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b154  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b155  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b156  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b157  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b158  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b159  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b128_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$4$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b16  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b160  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$5$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b161  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b162  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$5$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b163  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b164  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b165  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$5$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b166  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b167  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b168  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b169  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b17  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b170  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b171  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b172  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b173  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b174  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b175  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b176  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b177  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b178  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b179  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b18  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b180  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b181  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b182  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b183  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b184  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b185  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b186  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b187  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b188  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b189  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b19  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b190  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b191  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b160_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$5$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b192  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$6$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b193  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b194  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b195  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b196  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$6$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b197  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b198  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b199  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b2  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b20  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b200  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b201  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b202  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b203  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b204  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b205  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b206  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b207  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b208  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b209  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b21  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b210  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b211  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b212  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b213  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b214  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b215  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b216  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b217  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b218  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b219  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b22  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b220  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b221  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b222  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b223  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b192_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$6$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b224  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b225  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$7$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b226  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b227  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b228  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b229  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$7$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b23  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b230  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b231  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b232  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b233  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b234  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b235  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b236  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b237  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b238  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b239  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b24  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b240  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b241  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b242  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b243  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b244  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b245  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b246  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b247  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b248  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b249  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b25  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b250  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b251  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b252  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b253  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b254  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b255  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b224_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$7$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b256  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$8$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b257  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b258  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$8$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b259  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b26  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b260  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$8$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b261  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b262  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$8$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b263  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b264  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b265  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b266  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b267  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b268  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b269  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b27  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b270  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b271  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b272  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b273  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b274  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b275  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b276  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b277  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b278  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b279  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b28  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b280  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b281  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b282  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b283  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b284  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b285  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b286  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b287  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b256_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$8$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b288  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$9$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b289  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b29  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b290  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b291  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b292  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b293  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b294  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b295  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b296  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b297  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b298  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b299  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b3  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b30  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b300  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b301  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b302  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b303  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b304  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b305  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b306  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b307  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b308  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b309  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b31  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b310  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b311  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b312  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b313  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b314  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b315  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b316  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b317  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b318  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b319  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b288_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$9$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b32  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b320  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b321  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$10$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b322  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b323  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b324  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b325  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b326  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b327  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b328  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b329  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b33  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$1$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b330  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b331  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b332  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b333  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b334  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b335  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b336  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b337  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b338  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b339  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b34  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b340  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b341  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b342  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b343  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b344  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b345  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b346  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b347  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b348  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b349  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b35  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b350  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b351  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b320_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$10$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b352  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$11$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b353  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b354  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$11$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b355  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b356  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b357  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b358  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b359  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b36  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b360  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b361  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b362  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b363  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b364  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b365  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b366  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b367  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b368  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b369  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b37  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b370  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b371  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b372  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b373  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b374  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b375  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b376  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b377  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b378  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b379  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b38  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b380  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b381  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b382  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b383  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b352_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$11$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b384  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b385  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b386  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b387  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b388  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$12$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b389  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b39  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b390  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$12$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b391  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b392  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b393  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b394  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b395  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b396  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b397  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b398  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b399  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b4  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b40  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b400  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b401  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b402  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b403  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b404  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b405  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b406  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b407  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b408  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b409  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b41  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b410  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b411  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b412  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b413  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b414  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b415  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b384_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$12$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b416  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b417  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b418  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b419  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b42  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b420  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b421  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$13$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b422  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b423  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b424  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b425  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b426  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b427  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b428  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b429  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b43  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b430  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b431  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b432  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b433  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b434  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b435  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b436  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b437  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b438  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b439  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b44  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b440  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b441  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b442  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b443  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b444  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b445  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b446  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b447  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b416_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$13$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b448  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b449  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b45  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b450  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b451  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b452  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$14$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b453  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b454  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b455  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b456  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b457  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b458  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b459  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b46  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b460  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b461  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b462  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b463  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b464  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b465  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b466  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b467  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b468  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b469  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b47  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b470  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b471  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b472  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b473  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b474  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b475  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b476  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b477  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b478  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b479  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b448_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$14$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b48  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b480  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$15$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b481  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$15$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b482  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b483  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b484  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$15$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b485  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b486  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b487  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b488  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b489  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b49  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b490  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b491  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b492  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b493  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b494  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b495  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b496  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b497  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b498  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b499  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b5  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b50  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b500  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b501  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b502  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b503  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b504  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b505  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b506  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b507  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b508  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b509  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b51  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b510  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b511  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b480_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$15$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b512  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$16$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b513  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$16$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b514  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b515  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b516  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b517  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b518  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b519  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b52  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b520  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b521  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b522  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b523  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b524  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b525  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b526  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b527  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b528  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b529  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b53  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b530  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b531  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b532  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b533  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b534  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b535  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b536  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b537  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b538  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b539  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b54  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b540  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b541  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b542  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b543  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b512_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$16$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b544  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b545  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b546  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b547  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b548  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$17$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b549  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$17$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b55  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b550  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b551  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b552  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b553  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b554  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b555  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b556  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b557  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b558  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b559  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b56  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b560  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b561  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b562  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b563  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b564  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b565  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b566  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b567  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b568  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b569  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b57  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b570  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b571  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b572  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b573  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b574  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b575  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b544_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$17$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b576  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$18$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b577  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$18$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b578  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b579  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b58  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b580  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$18$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b581  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$18$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b582  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b583  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b584  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b585  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b586  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b587  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b588  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b589  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b59  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b590  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b591  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b592  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b593  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b594  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b595  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b596  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b597  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b598  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b599  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b6  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b60  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b600  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b601  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b602  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b603  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b604  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b605  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b606  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b607  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b576_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$18$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b608  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$19$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b609  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$19$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b61  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b610  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b611  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b612  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b613  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b614  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$19$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b615  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b616  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b617  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b618  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b619  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b62  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b620  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b621  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b622  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b623  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b624  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b625  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b626  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b627  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b628  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b629  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b63  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b32_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$1$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b630  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b631  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b632  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b633  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b634  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b635  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b636  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b637  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b638  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b639  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b608_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$19$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b64  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$2$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b640  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b641  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b642  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$20$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b643  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b644  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$20$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b645  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$20$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b646  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b647  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b648  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b649  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b65  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b650  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b651  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b652  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b653  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b654  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b655  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b656  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b657  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b658  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b659  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b66  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b660  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b661  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b662  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b663  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b664  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b665  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b666  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b667  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b668  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b669  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b67  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b670  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b671  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b640_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$20$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b672  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b673  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b674  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$21$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b675  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b676  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b677  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b678  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$21$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b679  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b68  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b680  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b681  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b682  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b683  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b684  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b685  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b686  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b687  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b688  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b689  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b69  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b690  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b691  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b692  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b693  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b694  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b695  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b696  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b697  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b698  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b699  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b7  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b70  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b700  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b701  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b702  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b703  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b672_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$21$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b704  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b705  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b706  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$22$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b707  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b708  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$22$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b709  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b71  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b710  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$22$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b711  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b712  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b713  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b714  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b715  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b716  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b717  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b718  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b719  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b72  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b720  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b721  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b722  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b723  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b724  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b725  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b726  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b727  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b728  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b729  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b73  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b730  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b731  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b732  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b733  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b734  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b735  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b704_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$22$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b736  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$23$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b737  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b738  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$23$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b739  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b74  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b740  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b741  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b742  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$23$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b743  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b744  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b745  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b746  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b747  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b748  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b749  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b75  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b750  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b751  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b752  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b753  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b754  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b755  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b756  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b757  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b758  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b759  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b76  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b760  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b761  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b762  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b763  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b764  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b765  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b766  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b767  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b736_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$23$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b768  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$24$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b769  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$24$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b77  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b770  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$24$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b771  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b772  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$24$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b773  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b774  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$24$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b775  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b776  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b777  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b778  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b779  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b78  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b780  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b781  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b782  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b783  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b784  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b785  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b786  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b787  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b788  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b789  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b79  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b790  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b791  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b792  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b793  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b794  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b795  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b796  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b797  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b798  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b799  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b768_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$24$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b8  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b80  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b800  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b801  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$25$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b802  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$25$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b803  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b804  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$25$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b805  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b806  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$25$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b807  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b808  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b809  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b81  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b810  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b811  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b812  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b813  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b814  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b815  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b816  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b817  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b818  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b819  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b82  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b820  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b821  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b822  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b823  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b824  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b825  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b826  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b827  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b828  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b829  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b83  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b830  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b831  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b800_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$25$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b832  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$26$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b833  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b834  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$26$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b835  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b836  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b837  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$26$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b838  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$26$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b839  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b84  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b840  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b841  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b842  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b843  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b844  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b845  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b846  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b847  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b848  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b849  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b85  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b850  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b851  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b852  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b853  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b854  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b855  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b856  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b857  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b858  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b859  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b86  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b860  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b861  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b862  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b863  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b832_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$26$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b864  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b865  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$27$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b866  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$27$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b867  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b868  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b869  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$27$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b87  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b870  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$27$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b871  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b872  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b873  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b874  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b875  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b876  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b877  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b878  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b879  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b88  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b880  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b881  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b882  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b883  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b884  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b885  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b886  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b887  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b888  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b889  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b89  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b890  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b891  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b892  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b893  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b894  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b895  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b864_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$27$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b896  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b897  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$28$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b898  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b899  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b9  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b0_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$0$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b90  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b900  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$28$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b901  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b902  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b903  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b904  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b905  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b906  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b907  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b908  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b909  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b91  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b910  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b911  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b912  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b913  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b914  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b915  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b916  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b917  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b918  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b919  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b92  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b920  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b921  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b922  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b923  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b924  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b925  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b926  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b927  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b896_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$28$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b928  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$29$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b929  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b93  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b930  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$29$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b931  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b932  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$29$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b933  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$29$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b934  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$29$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b935  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b936  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b937  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b938  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b939  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b94  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b940  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b941  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b942  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b943  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b944  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b945  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b946  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b947  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b948  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b949  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b95  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b64_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$2$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b950  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b951  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b952  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b953  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b954  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b955  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b956  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b957  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b958  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b959  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b928_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$29$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b96  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b960  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$30$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b961  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$30$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b962  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$30$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b963  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b964  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$30$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b965  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$30$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b966  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$30$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b967  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [7]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b968  (
    .clk(clock),
    .d(\t/a/reg_writedat [8]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [8]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b969  (
    .clk(clock),
    .d(\t/a/reg_writedat [9]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [9]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b97  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b970  (
    .clk(clock),
    .d(\t/a/reg_writedat [10]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [10]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b971  (
    .clk(clock),
    .d(\t/a/reg_writedat [11]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [11]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b972  (
    .clk(clock),
    .d(\t/a/reg_writedat [12]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [12]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b973  (
    .clk(clock),
    .d(\t/a/reg_writedat [13]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [13]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b974  (
    .clk(clock),
    .d(\t/a/reg_writedat [14]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [14]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b975  (
    .clk(clock),
    .d(\t/a/reg_writedat [15]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [15]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b976  (
    .clk(clock),
    .d(\t/a/reg_writedat [16]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [16]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b977  (
    .clk(clock),
    .d(\t/a/reg_writedat [17]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [17]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b978  (
    .clk(clock),
    .d(\t/a/reg_writedat [18]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [18]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b979  (
    .clk(clock),
    .d(\t/a/reg_writedat [19]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [19]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b98  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b980  (
    .clk(clock),
    .d(\t/a/reg_writedat [20]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [20]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b981  (
    .clk(clock),
    .d(\t/a/reg_writedat [21]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [21]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b982  (
    .clk(clock),
    .d(\t/a/reg_writedat [22]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [22]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b983  (
    .clk(clock),
    .d(\t/a/reg_writedat [23]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [23]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b984  (
    .clk(clock),
    .d(\t/a/reg_writedat [24]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [24]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b985  (
    .clk(clock),
    .d(\t/a/reg_writedat [25]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [25]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b986  (
    .clk(clock),
    .d(\t/a/reg_writedat [26]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [26]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b987  (
    .clk(clock),
    .d(\t/a/reg_writedat [27]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [27]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b988  (
    .clk(clock),
    .d(\t/a/reg_writedat [28]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [28]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b989  (
    .clk(clock),
    .d(\t/a/reg_writedat [29]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [29]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b99  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b100_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$3$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b990  (
    .clk(clock),
    .d(\t/a/reg_writedat [30]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [30]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b991  (
    .clk(clock),
    .d(\t/a/reg_writedat [31]),
    .en(\t/a/regfile/mux39_b960_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$30$ [31]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b992  (
    .clk(clock),
    .d(\t/a/reg_writedat [0]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$31$ [0]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b993  (
    .clk(clock),
    .d(\t/a/reg_writedat [1]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$31$ [1]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b994  (
    .clk(clock),
    .d(\t/a/reg_writedat [2]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$31$ [2]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b995  (
    .clk(clock),
    .d(\t/a/reg_writedat [3]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [3]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b996  (
    .clk(clock),
    .d(\t/a/reg_writedat [4]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [4]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b997  (
    .clk(clock),
    .d(\t/a/reg_writedat [5]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(1'b0),
    .set(~rst),
    .q(\t/a/regfile/regfile$31$ [5]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b998  (
    .clk(clock),
    .d(\t/a/reg_writedat [6]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [6]));  // register.v(63)
  reg_ar_as_w1 \t/a/regfile/reg0_b999  (
    .clk(clock),
    .d(\t/a/reg_writedat [7]),
    .en(\t/a/regfile/mux39_b1000_sel_is_3_o ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/a/regfile/regfile$31$ [7]));  // register.v(63)
  not \t/a/regfile/u10  (\t/a/regfile/n40 , \t/a/WB_rd [2]);  // register.v(63)
  and \t/a/regfile/u11  (\t/a/regfile/n6 , \t/a/regfile/n0 , \t/a/regfile/n3 );  // register.v(18)
  and \t/a/regfile/u12  (\t/a/regfile/n30 , \t/a/regfile/n33 , \t/a/WB_rd [2]);  // register.v(63)
  and \t/a/regfile/u13  (\t/a/regfile/n31 , \t/a/regfile/n35 , \t/a/regfile/n40 );  // register.v(63)
  not \t/a/regfile/u14  (\t/a/regfile/n80 , \t/a/WB_rd [1]);  // register.v(63)
  and \t/a/regfile/u15  (\t/a/regfile/n34 , \t/a/WB_rd [0], \t/a/WB_rd [1]);  // register.v(63)
  not \t/a/regfile/u17  (\t/a/regfile/n37 , \t/a/WB_rd [0]);  // register.v(63)
  and \t/a/regfile/u18  (\t/a/regfile/n29 , \t/a/regfile/n33 , \t/a/regfile/n40 );  // register.v(63)
  and \t/a/regfile/u19  (\t/a/regfile/n28 , \t/a/regfile/n36 , \t/a/WB_rd [2]);  // register.v(63)
  and \t/a/regfile/u2  (\t/a/regfile/n32 , \t/a/regfile/n35 , \t/a/WB_rd [2]);  // register.v(63)
  and \t/a/regfile/u20  (\t/a/regfile/n27 , \t/a/regfile/n36 , \t/a/regfile/n40 );  // register.v(63)
  and \t/a/regfile/u21  (\t/a/regfile/n26 , \t/a/regfile/n34 , \t/a/WB_rd [2]);  // register.v(63)
  and \t/a/regfile/u22  (\t/a/regfile/n25 , \t/a/regfile/n34 , \t/a/regfile/n40 );  // register.v(63)
  and \t/a/regfile/u23  (\t/a/regfile/n24 , \t/a/regfile/n31 , \t/a/WB_rd [3]);  // register.v(63)
  and \t/a/regfile/u24  (\t/a/regfile/n23 , \t/a/regfile/n31 , \t/a/regfile/n39 );  // register.v(63)
  and \t/a/regfile/u25  (\t/a/regfile/n22 , \t/a/regfile/n29 , \t/a/WB_rd [3]);  // register.v(63)
  and \t/a/regfile/u26  (\t/a/regfile/n21 , \t/a/regfile/n29 , \t/a/regfile/n39 );  // register.v(63)
  and \t/a/regfile/u27  (\t/a/regfile/n20 , \t/a/regfile/n27 , \t/a/WB_rd [3]);  // register.v(63)
  and \t/a/regfile/u28  (\t/a/regfile/n19 , \t/a/regfile/n27 , \t/a/regfile/n39 );  // register.v(63)
  and \t/a/regfile/u29  (\t/a/regfile/n18 , \t/a/regfile/n25 , \t/a/WB_rd [3]);  // register.v(63)
  and \t/a/regfile/u3  (\t/a/regfile/n33 , \t/a/WB_rd [0], \t/a/regfile/n80 );  // register.v(63)
  and \t/a/regfile/u30  (\t/a/regfile/n17 , \t/a/regfile/n25 , \t/a/regfile/n39 );  // register.v(63)
  and \t/a/regfile/u31  (\t/a/regfile/n16 , \t/a/regfile/n32 , \t/a/WB_rd [3]);  // register.v(63)
  and \t/a/regfile/u32  (\t/a/regfile/n15 , \t/a/regfile/n32 , \t/a/regfile/n39 );  // register.v(63)
  and \t/a/regfile/u33  (\t/a/regfile/n14 , \t/a/regfile/n30 , \t/a/WB_rd [3]);  // register.v(63)
  and \t/a/regfile/u34  (\t/a/regfile/n13 , \t/a/regfile/n30 , \t/a/regfile/n39 );  // register.v(63)
  and \t/a/regfile/u35  (\t/a/regfile/n12 , \t/a/regfile/n28 , \t/a/WB_rd [3]);  // register.v(63)
  and \t/a/regfile/u36  (\t/a/regfile/n11 , \t/a/regfile/n28 , \t/a/regfile/n39 );  // register.v(63)
  and \t/a/regfile/u37  (\t/a/regfile/n10 , \t/a/regfile/n26 , \t/a/WB_rd [3]);  // register.v(63)
  and \t/a/regfile/u38  (\t/a/regfile/n9 , \t/a/regfile/n26 , \t/a/regfile/n39 );  // register.v(63)
  and \t/a/regfile/u39  (\t/a/regfile/n46 [16], \t/a/regfile/n23 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u4  (\t/a/regfile/n2 , \t/a/regfile/n0 , \t/a/regfile/n1 );  // register.v(10)
  and \t/a/regfile/u40  (\t/a/regfile/n46 [0], \t/a/regfile/n23 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u41  (\t/a/regfile/n46 [17], \t/a/regfile/n21 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u42  (\t/a/regfile/n46 [1], \t/a/regfile/n21 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u43  (\t/a/regfile/n46 [18], \t/a/regfile/n19 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u44  (\t/a/regfile/n46 [2], \t/a/regfile/n19 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u45  (\t/a/regfile/n46 [19], \t/a/regfile/n17 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u46  (\t/a/regfile/n46 [3], \t/a/regfile/n17 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u47  (\t/a/regfile/n46 [20], \t/a/regfile/n15 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u48  (\t/a/regfile/n46 [4], \t/a/regfile/n15 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u49  (\t/a/regfile/n46 [21], \t/a/regfile/n13 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u5  (\t/a/regfile/n4 , \t/a/regfile/n2 , \t/a/regfile/n3 );  // register.v(10)
  and \t/a/regfile/u50  (\t/a/regfile/n46 [5], \t/a/regfile/n13 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u51  (\t/a/regfile/n46 [22], \t/a/regfile/n11 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u52  (\t/a/regfile/n46 [6], \t/a/regfile/n11 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u53  (\t/a/regfile/n46 [23], \t/a/regfile/n9 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u54  (\t/a/regfile/n46 [7], \t/a/regfile/n9 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u55  (\t/a/regfile/n46 [24], \t/a/regfile/n24 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u56  (\t/a/regfile/n46 [8], \t/a/regfile/n24 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u57  (\t/a/regfile/n46 [25], \t/a/regfile/n22 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u58  (\t/a/regfile/n46 [9], \t/a/regfile/n22 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u59  (\t/a/regfile/n46 [26], \t/a/regfile/n20 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u6  (\t/a/regfile/n35 , \t/a/regfile/n37 , \t/a/regfile/n80 );  // register.v(63)
  and \t/a/regfile/u60  (\t/a/regfile/n46 [10], \t/a/regfile/n20 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u61  (\t/a/regfile/n46 [27], \t/a/regfile/n18 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u62  (\t/a/regfile/n46 [11], \t/a/regfile/n18 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u63  (\t/a/regfile/n46 [28], \t/a/regfile/n16 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u64  (\t/a/regfile/n46 [12], \t/a/regfile/n16 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u65  (\t/a/regfile/n46 [29], \t/a/regfile/n14 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u66  (\t/a/regfile/n46 [13], \t/a/regfile/n14 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u67  (\t/a/regfile/n46 [30], \t/a/regfile/n12 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u68  (\t/a/regfile/n46 [14], \t/a/regfile/n12 , \t/a/regfile/n38 );  // register.v(63)
  and \t/a/regfile/u69  (\t/a/regfile/n46 [31], \t/a/regfile/n10 , \t/a/WB_rd [4]);  // register.v(63)
  and \t/a/regfile/u7  (\t/a/regfile/n36 , \t/a/regfile/n37 , \t/a/WB_rd [1]);  // register.v(63)
  and \t/a/regfile/u70  (\t/a/regfile/n46 [15], \t/a/regfile/n10 , \t/a/regfile/n38 );  // register.v(63)
  not \t/a/regfile/u8  (\t/a/regfile/n38 , \t/a/WB_rd [4]);  // register.v(63)
  not \t/a/regfile/u9  (\t/a/regfile/n39 , \t/a/WB_rd [3]);  // register.v(63)
  eq_w1 \t/a/risk_jump/eq1  (
    .i0(\t/a/risk_jump/EX_risk ),
    .i1(1'b1),
    .o(\t/a/risk_jump/n10 ));  // PC.v(176)
  eq_w5 \t/a/risk_jump/eq2  (
    .i0(\t/a/EX_rd ),
    .i1(\t/a/ID_rs1 ),
    .o(\t/a/risk_jump/n11 ));  // PC.v(177)
  eq_w1 \t/a/risk_jump/eq3  (
    .i0(\t/a/risk_jump/MEM_risk ),
    .i1(1'b1),
    .o(\t/a/risk_jump/n17 ));  // PC.v(181)
  eq_w5 \t/a/risk_jump/eq4  (
    .i0(\t/a/MEM_rd ),
    .i1(\t/a/ID_rs1 ),
    .o(\t/a/risk_jump/n24 ));  // PC.v(185)
  eq_w1 \t/a/risk_jump/eq5  (
    .i0(\t/a/risk_jump/WB_risk ),
    .i1(1'b1),
    .o(\t/a/risk_jump/n26 ));  // PC.v(187)
  eq_w5 \t/a/risk_jump/eq7  (
    .i0(\t/a/EX_rd ),
    .i1(\t/a/ID_rs2 ),
    .o(\t/a/risk_jump/n35 ));  // PC.v(208)
  eq_w5 \t/a/risk_jump/eq8  (
    .i0(\t/a/MEM_rd ),
    .i1(\t/a/ID_rs2 ),
    .o(\t/a/risk_jump/n42 ));  // PC.v(216)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b0  (
    .i0(\t/a/ID_read_dat1 [0]),
    .i1(\t/a/aludat [0]),
    .i2(\t/a/MEM_aludat [0]),
    .i3(\t/a/reg_writedat [0]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [0]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b1  (
    .i0(\t/a/ID_read_dat1 [1]),
    .i1(\t/a/aludat [1]),
    .i2(\t/a/MEM_aludat [1]),
    .i3(\t/a/reg_writedat [1]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [1]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b10  (
    .i0(\t/a/ID_read_dat1 [10]),
    .i1(\t/a/aludat [10]),
    .i2(\t/a/MEM_aludat [10]),
    .i3(\t/a/reg_writedat [10]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [10]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b11  (
    .i0(\t/a/ID_read_dat1 [11]),
    .i1(\t/a/aludat [11]),
    .i2(\t/a/MEM_aludat [11]),
    .i3(\t/a/reg_writedat [11]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [11]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b12  (
    .i0(\t/a/ID_read_dat1 [12]),
    .i1(\t/a/aludat [12]),
    .i2(\t/a/MEM_aludat [12]),
    .i3(\t/a/reg_writedat [12]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [12]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b13  (
    .i0(\t/a/ID_read_dat1 [13]),
    .i1(\t/a/aludat [13]),
    .i2(\t/a/MEM_aludat [13]),
    .i3(\t/a/reg_writedat [13]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [13]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b14  (
    .i0(\t/a/ID_read_dat1 [14]),
    .i1(\t/a/aludat [14]),
    .i2(\t/a/MEM_aludat [14]),
    .i3(\t/a/reg_writedat [14]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [14]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b15  (
    .i0(\t/a/ID_read_dat1 [15]),
    .i1(\t/a/aludat [15]),
    .i2(\t/a/MEM_aludat [15]),
    .i3(\t/a/reg_writedat [15]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [15]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b16  (
    .i0(\t/a/ID_read_dat1 [16]),
    .i1(\t/a/aludat [16]),
    .i2(\t/a/MEM_aludat [16]),
    .i3(\t/a/reg_writedat [16]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [16]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b17  (
    .i0(\t/a/ID_read_dat1 [17]),
    .i1(\t/a/aludat [17]),
    .i2(\t/a/MEM_aludat [17]),
    .i3(\t/a/reg_writedat [17]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [17]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b18  (
    .i0(\t/a/ID_read_dat1 [18]),
    .i1(\t/a/aludat [18]),
    .i2(\t/a/MEM_aludat [18]),
    .i3(\t/a/reg_writedat [18]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [18]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b19  (
    .i0(\t/a/ID_read_dat1 [19]),
    .i1(\t/a/aludat [19]),
    .i2(\t/a/MEM_aludat [19]),
    .i3(\t/a/reg_writedat [19]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [19]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b2  (
    .i0(\t/a/ID_read_dat1 [2]),
    .i1(\t/a/aludat [2]),
    .i2(\t/a/MEM_aludat [2]),
    .i3(\t/a/reg_writedat [2]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [2]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b20  (
    .i0(\t/a/ID_read_dat1 [20]),
    .i1(\t/a/aludat [20]),
    .i2(\t/a/MEM_aludat [20]),
    .i3(\t/a/reg_writedat [20]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [20]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b21  (
    .i0(\t/a/ID_read_dat1 [21]),
    .i1(\t/a/aludat [21]),
    .i2(\t/a/MEM_aludat [21]),
    .i3(\t/a/reg_writedat [21]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [21]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b22  (
    .i0(\t/a/ID_read_dat1 [22]),
    .i1(\t/a/aludat [22]),
    .i2(\t/a/MEM_aludat [22]),
    .i3(\t/a/reg_writedat [22]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [22]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b23  (
    .i0(\t/a/ID_read_dat1 [23]),
    .i1(\t/a/aludat [23]),
    .i2(\t/a/MEM_aludat [23]),
    .i3(\t/a/reg_writedat [23]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [23]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b24  (
    .i0(\t/a/ID_read_dat1 [24]),
    .i1(\t/a/aludat [24]),
    .i2(\t/a/MEM_aludat [24]),
    .i3(\t/a/reg_writedat [24]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [24]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b25  (
    .i0(\t/a/ID_read_dat1 [25]),
    .i1(\t/a/aludat [25]),
    .i2(\t/a/MEM_aludat [25]),
    .i3(\t/a/reg_writedat [25]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [25]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b26  (
    .i0(\t/a/ID_read_dat1 [26]),
    .i1(\t/a/aludat [26]),
    .i2(\t/a/MEM_aludat [26]),
    .i3(\t/a/reg_writedat [26]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [26]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b27  (
    .i0(\t/a/ID_read_dat1 [27]),
    .i1(\t/a/aludat [27]),
    .i2(\t/a/MEM_aludat [27]),
    .i3(\t/a/reg_writedat [27]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [27]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b28  (
    .i0(\t/a/ID_read_dat1 [28]),
    .i1(\t/a/aludat [28]),
    .i2(\t/a/MEM_aludat [28]),
    .i3(\t/a/reg_writedat [28]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [28]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b29  (
    .i0(\t/a/ID_read_dat1 [29]),
    .i1(\t/a/aludat [29]),
    .i2(\t/a/MEM_aludat [29]),
    .i3(\t/a/reg_writedat [29]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [29]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b3  (
    .i0(\t/a/ID_read_dat1 [3]),
    .i1(\t/a/aludat [3]),
    .i2(\t/a/MEM_aludat [3]),
    .i3(\t/a/reg_writedat [3]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [3]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b30  (
    .i0(\t/a/ID_read_dat1 [30]),
    .i1(\t/a/aludat [30]),
    .i2(\t/a/MEM_aludat [30]),
    .i3(\t/a/reg_writedat [30]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [30]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b31  (
    .i0(\t/a/ID_read_dat1 [31]),
    .i1(\t/a/aludat [31]),
    .i2(\t/a/MEM_aludat [31]),
    .i3(\t/a/reg_writedat [31]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [31]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b4  (
    .i0(\t/a/ID_read_dat1 [4]),
    .i1(\t/a/aludat [4]),
    .i2(\t/a/MEM_aludat [4]),
    .i3(\t/a/reg_writedat [4]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [4]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b5  (
    .i0(\t/a/ID_read_dat1 [5]),
    .i1(\t/a/aludat [5]),
    .i2(\t/a/MEM_aludat [5]),
    .i3(\t/a/reg_writedat [5]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [5]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b6  (
    .i0(\t/a/ID_read_dat1 [6]),
    .i1(\t/a/aludat [6]),
    .i2(\t/a/MEM_aludat [6]),
    .i3(\t/a/reg_writedat [6]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [6]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b7  (
    .i0(\t/a/ID_read_dat1 [7]),
    .i1(\t/a/aludat [7]),
    .i2(\t/a/MEM_aludat [7]),
    .i3(\t/a/reg_writedat [7]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [7]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b8  (
    .i0(\t/a/ID_read_dat1 [8]),
    .i1(\t/a/aludat [8]),
    .i2(\t/a/MEM_aludat [8]),
    .i3(\t/a/reg_writedat [8]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [8]));  // PC.v(172)
  binary_mux_s2_w1 \t/a/risk_jump/mux0_b9  (
    .i0(\t/a/ID_read_dat1 [9]),
    .i1(\t/a/aludat [9]),
    .i2(\t/a/MEM_aludat [9]),
    .i3(\t/a/reg_writedat [9]),
    .sel(\t/a/risk_jump/rs1_select ),
    .o(\t/a/ID_jump_regdat1 [9]));  // PC.v(172)
  binary_mux_s1_w1 \t/a/risk_jump/mux1_b0  (
    .i0(\t/a/risk_jump/n33 ),
    .i1(1'b0),
    .sel(\t/a/risk_jump/n25 ),
    .o(\t/a/risk_jump/n34 [0]));  // PC.v(194)
  binary_mux_s1_w1 \t/a/risk_jump/mux1_b1  (
    .i0(\t/a/risk_jump/n33 ),
    .i1(1'b1),
    .sel(\t/a/risk_jump/n25 ),
    .o(\t/a/risk_jump/n34 [1]));  // PC.v(194)
  binary_mux_s1_w1 \t/a/risk_jump/mux2_b0  (
    .i0(\t/a/risk_jump/n34 [0]),
    .i1(1'b1),
    .sel(\t/a/risk_jump/n16 ),
    .o(\t/a/risk_jump/rs1_select [0]));  // PC.v(194)
  binary_mux_s1_w1 \t/a/risk_jump/mux2_b1  (
    .i0(\t/a/risk_jump/n34 [1]),
    .i1(1'b0),
    .sel(\t/a/risk_jump/n16 ),
    .o(\t/a/risk_jump/rs1_select [1]));  // PC.v(194)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b0  (
    .i0(\t/a/ID_read_dat2 [0]),
    .i1(\t/a/aludat [0]),
    .i2(\t/a/MEM_aludat [0]),
    .i3(\t/a/reg_writedat [0]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [0]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b1  (
    .i0(\t/a/ID_read_dat2 [1]),
    .i1(\t/a/aludat [1]),
    .i2(\t/a/MEM_aludat [1]),
    .i3(\t/a/reg_writedat [1]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [1]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b10  (
    .i0(\t/a/ID_read_dat2 [10]),
    .i1(\t/a/aludat [10]),
    .i2(\t/a/MEM_aludat [10]),
    .i3(\t/a/reg_writedat [10]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [10]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b11  (
    .i0(\t/a/ID_read_dat2 [11]),
    .i1(\t/a/aludat [11]),
    .i2(\t/a/MEM_aludat [11]),
    .i3(\t/a/reg_writedat [11]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [11]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b12  (
    .i0(\t/a/ID_read_dat2 [12]),
    .i1(\t/a/aludat [12]),
    .i2(\t/a/MEM_aludat [12]),
    .i3(\t/a/reg_writedat [12]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [12]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b13  (
    .i0(\t/a/ID_read_dat2 [13]),
    .i1(\t/a/aludat [13]),
    .i2(\t/a/MEM_aludat [13]),
    .i3(\t/a/reg_writedat [13]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [13]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b14  (
    .i0(\t/a/ID_read_dat2 [14]),
    .i1(\t/a/aludat [14]),
    .i2(\t/a/MEM_aludat [14]),
    .i3(\t/a/reg_writedat [14]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [14]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b15  (
    .i0(\t/a/ID_read_dat2 [15]),
    .i1(\t/a/aludat [15]),
    .i2(\t/a/MEM_aludat [15]),
    .i3(\t/a/reg_writedat [15]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [15]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b16  (
    .i0(\t/a/ID_read_dat2 [16]),
    .i1(\t/a/aludat [16]),
    .i2(\t/a/MEM_aludat [16]),
    .i3(\t/a/reg_writedat [16]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [16]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b17  (
    .i0(\t/a/ID_read_dat2 [17]),
    .i1(\t/a/aludat [17]),
    .i2(\t/a/MEM_aludat [17]),
    .i3(\t/a/reg_writedat [17]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [17]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b18  (
    .i0(\t/a/ID_read_dat2 [18]),
    .i1(\t/a/aludat [18]),
    .i2(\t/a/MEM_aludat [18]),
    .i3(\t/a/reg_writedat [18]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [18]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b19  (
    .i0(\t/a/ID_read_dat2 [19]),
    .i1(\t/a/aludat [19]),
    .i2(\t/a/MEM_aludat [19]),
    .i3(\t/a/reg_writedat [19]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [19]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b2  (
    .i0(\t/a/ID_read_dat2 [2]),
    .i1(\t/a/aludat [2]),
    .i2(\t/a/MEM_aludat [2]),
    .i3(\t/a/reg_writedat [2]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [2]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b20  (
    .i0(\t/a/ID_read_dat2 [20]),
    .i1(\t/a/aludat [20]),
    .i2(\t/a/MEM_aludat [20]),
    .i3(\t/a/reg_writedat [20]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [20]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b21  (
    .i0(\t/a/ID_read_dat2 [21]),
    .i1(\t/a/aludat [21]),
    .i2(\t/a/MEM_aludat [21]),
    .i3(\t/a/reg_writedat [21]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [21]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b22  (
    .i0(\t/a/ID_read_dat2 [22]),
    .i1(\t/a/aludat [22]),
    .i2(\t/a/MEM_aludat [22]),
    .i3(\t/a/reg_writedat [22]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [22]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b23  (
    .i0(\t/a/ID_read_dat2 [23]),
    .i1(\t/a/aludat [23]),
    .i2(\t/a/MEM_aludat [23]),
    .i3(\t/a/reg_writedat [23]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [23]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b24  (
    .i0(\t/a/ID_read_dat2 [24]),
    .i1(\t/a/aludat [24]),
    .i2(\t/a/MEM_aludat [24]),
    .i3(\t/a/reg_writedat [24]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [24]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b25  (
    .i0(\t/a/ID_read_dat2 [25]),
    .i1(\t/a/aludat [25]),
    .i2(\t/a/MEM_aludat [25]),
    .i3(\t/a/reg_writedat [25]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [25]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b26  (
    .i0(\t/a/ID_read_dat2 [26]),
    .i1(\t/a/aludat [26]),
    .i2(\t/a/MEM_aludat [26]),
    .i3(\t/a/reg_writedat [26]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [26]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b27  (
    .i0(\t/a/ID_read_dat2 [27]),
    .i1(\t/a/aludat [27]),
    .i2(\t/a/MEM_aludat [27]),
    .i3(\t/a/reg_writedat [27]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [27]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b28  (
    .i0(\t/a/ID_read_dat2 [28]),
    .i1(\t/a/aludat [28]),
    .i2(\t/a/MEM_aludat [28]),
    .i3(\t/a/reg_writedat [28]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [28]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b29  (
    .i0(\t/a/ID_read_dat2 [29]),
    .i1(\t/a/aludat [29]),
    .i2(\t/a/MEM_aludat [29]),
    .i3(\t/a/reg_writedat [29]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [29]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b3  (
    .i0(\t/a/ID_read_dat2 [3]),
    .i1(\t/a/aludat [3]),
    .i2(\t/a/MEM_aludat [3]),
    .i3(\t/a/reg_writedat [3]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [3]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b30  (
    .i0(\t/a/ID_read_dat2 [30]),
    .i1(\t/a/aludat [30]),
    .i2(\t/a/MEM_aludat [30]),
    .i3(\t/a/reg_writedat [30]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [30]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b31  (
    .i0(\t/a/ID_read_dat2 [31]),
    .i1(\t/a/aludat [31]),
    .i2(\t/a/MEM_aludat [31]),
    .i3(\t/a/reg_writedat [31]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [31]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b4  (
    .i0(\t/a/ID_read_dat2 [4]),
    .i1(\t/a/aludat [4]),
    .i2(\t/a/MEM_aludat [4]),
    .i3(\t/a/reg_writedat [4]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [4]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b5  (
    .i0(\t/a/ID_read_dat2 [5]),
    .i1(\t/a/aludat [5]),
    .i2(\t/a/MEM_aludat [5]),
    .i3(\t/a/reg_writedat [5]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [5]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b6  (
    .i0(\t/a/ID_read_dat2 [6]),
    .i1(\t/a/aludat [6]),
    .i2(\t/a/MEM_aludat [6]),
    .i3(\t/a/reg_writedat [6]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [6]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b7  (
    .i0(\t/a/ID_read_dat2 [7]),
    .i1(\t/a/aludat [7]),
    .i2(\t/a/MEM_aludat [7]),
    .i3(\t/a/reg_writedat [7]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [7]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b8  (
    .i0(\t/a/ID_read_dat2 [8]),
    .i1(\t/a/aludat [8]),
    .i2(\t/a/MEM_aludat [8]),
    .i3(\t/a/reg_writedat [8]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [8]));  // PC.v(203)
  binary_mux_s2_w1 \t/a/risk_jump/mux3_b9  (
    .i0(\t/a/ID_read_dat2 [9]),
    .i1(\t/a/aludat [9]),
    .i2(\t/a/MEM_aludat [9]),
    .i3(\t/a/reg_writedat [9]),
    .sel(\t/a/risk_jump/rs2_select ),
    .o(\t/a/ID_jump_regdat2 [9]));  // PC.v(203)
  binary_mux_s1_w1 \t/a/risk_jump/mux4_b0  (
    .i0(\t/a/risk_jump/n48 ),
    .i1(1'b0),
    .sel(\t/a/risk_jump/n43 ),
    .o(\t/a/risk_jump/n49 [0]));  // PC.v(225)
  binary_mux_s1_w1 \t/a/risk_jump/mux4_b1  (
    .i0(\t/a/risk_jump/n48 ),
    .i1(1'b1),
    .sel(\t/a/risk_jump/n43 ),
    .o(\t/a/risk_jump/n49 [1]));  // PC.v(225)
  binary_mux_s1_w1 \t/a/risk_jump/mux5_b0  (
    .i0(\t/a/risk_jump/n49 [0]),
    .i1(1'b1),
    .sel(\t/a/risk_jump/n38 ),
    .o(\t/a/risk_jump/rs2_select [0]));  // PC.v(225)
  binary_mux_s1_w1 \t/a/risk_jump/mux5_b1  (
    .i0(\t/a/risk_jump/n49 [1]),
    .i1(1'b0),
    .sel(\t/a/risk_jump/n38 ),
    .o(\t/a/risk_jump/rs2_select [1]));  // PC.v(225)
  ne_w7 \t/a/risk_jump/neq0  (
    .i0(\t/a/EX_op ),
    .i1(7'b0100011),
    .o(\t/a/risk_jump/n1 ));  // PC.v(143)
  ne_w7 \t/a/risk_jump/neq1  (
    .i0(\t/a/EX_op ),
    .i1(7'b1100011),
    .o(\t/a/risk_jump/n3 ));  // PC.v(144)
  ne_w5 \t/a/risk_jump/neq12  (
    .i0(\t/a/MEM_rd ),
    .i1(\t/a/ID_rs1 ),
    .o(\t/a/risk_jump/n30 ));  // PC.v(190)
  ne_w5 \t/a/risk_jump/neq13  (
    .i0(\t/a/EX_rd ),
    .i1(\t/a/ID_rs2 ),
    .o(\t/a/risk_jump/n39 ));  // PC.v(214)
  ne_w5 \t/a/risk_jump/neq14  (
    .i0(\t/a/MEM_rd ),
    .i1(\t/a/ID_rs2 ),
    .o(\t/a/risk_jump/n45 ));  // PC.v(221)
  ne_w5 \t/a/risk_jump/neq6  (
    .i0(\t/a/EX_rd ),
    .i1(5'b00000),
    .o(\t/a/risk_jump/n13 ));  // PC.v(178)
  ne_w7 \t/a/risk_jump/neq7  (
    .i0(\t/a/EX_op ),
    .i1(7'b0000011),
    .o(\t/a/risk_jump/n15 ));  // PC.v(179)
  ne_w5 \t/a/risk_jump/neq9  (
    .i0(\t/a/EX_rd ),
    .i1(\t/a/ID_rs1 ),
    .o(\t/a/risk_jump/n20 ));  // PC.v(183)
  and \t/a/risk_jump/u10  (\t/a/risk_jump/n16 , \t/a/risk_jump/n14 , \t/a/risk_jump/n15 );  // PC.v(179)
  and \t/a/risk_jump/u11  (\t/a/risk_jump/n19 , \t/a/risk_jump/n17 , \t/a/n11 );  // PC.v(182)
  and \t/a/risk_jump/u12  (\t/a/risk_jump/n21 , \t/a/risk_jump/n19 , \t/a/risk_jump/n20 );  // PC.v(183)
  and \t/a/risk_jump/u13  (\t/a/risk_jump/n23 , \t/a/risk_jump/n21 , \t/a/n13 );  // PC.v(184)
  and \t/a/risk_jump/u14  (\t/a/risk_jump/n25 , \t/a/risk_jump/n23 , \t/a/risk_jump/n24 );  // PC.v(185)
  and \t/a/risk_jump/u15  (\t/a/risk_jump/n28 , \t/a/risk_jump/n26 , \t/a/n18 );  // PC.v(188)
  and \t/a/risk_jump/u16  (\t/a/risk_jump/n29 , \t/a/risk_jump/n28 , \t/a/risk_jump/n20 );  // PC.v(189)
  and \t/a/risk_jump/u17  (\t/a/risk_jump/n31 , \t/a/risk_jump/n29 , \t/a/risk_jump/n30 );  // PC.v(190)
  and \t/a/risk_jump/u18  (\t/a/risk_jump/n33 , \t/a/risk_jump/n31 , \t/a/regfile/n1 );  // PC.v(192)
  and \t/a/risk_jump/u19  (\t/a/risk_jump/n36 , \t/a/risk_jump/n10 , \t/a/risk_jump/n35 );  // PC.v(208)
  and \t/a/risk_jump/u2  (\t/a/risk_jump/n2 , \t/a/condition/n1 , \t/a/risk_jump/n1 );  // PC.v(143)
  and \t/a/risk_jump/u20  (\t/a/risk_jump/n37 , \t/a/risk_jump/n36 , \t/a/risk_jump/n13 );  // PC.v(209)
  and \t/a/risk_jump/u21  (\t/a/risk_jump/n38 , \t/a/risk_jump/n37 , \t/a/risk_jump/n15 );  // PC.v(210)
  and \t/a/risk_jump/u22  (\t/a/risk_jump/n40 , \t/a/risk_jump/n19 , \t/a/risk_jump/n39 );  // PC.v(214)
  and \t/a/risk_jump/u23  (\t/a/risk_jump/n41 , \t/a/risk_jump/n40 , \t/a/n13 );  // PC.v(215)
  and \t/a/risk_jump/u24  (\t/a/risk_jump/n43 , \t/a/risk_jump/n41 , \t/a/risk_jump/n42 );  // PC.v(216)
  and \t/a/risk_jump/u25  (\t/a/risk_jump/n44 , \t/a/risk_jump/n28 , \t/a/risk_jump/n39 );  // PC.v(220)
  and \t/a/risk_jump/u26  (\t/a/risk_jump/n46 , \t/a/risk_jump/n44 , \t/a/risk_jump/n45 );  // PC.v(221)
  and \t/a/risk_jump/u27  (\t/a/risk_jump/n48 , \t/a/risk_jump/n46 , \t/a/regfile/n3 );  // PC.v(223)
  and \t/a/risk_jump/u28  (\t/a/risk_jump/n51 , \t/a/condition/n1 , \t/a/aluin/n11 );  // PC.v(230)
  or \t/a/risk_jump/u29  (\t/a/risk_jump/n52 , \t/a/risk_jump/n11 , \t/a/risk_jump/n35 );  // PC.v(232)
  and \t/a/risk_jump/u3  (\t/a/risk_jump/EX_risk , \t/a/risk_jump/n2 , \t/a/risk_jump/n3 );  // PC.v(144)
  and \t/a/risk_jump/u30  (\t/a/risk_jump/n53 , \t/a/risk_jump/n51 , \t/a/risk_jump/n52 );  // PC.v(232)
  and \t/a/risk_jump/u31  (\t/a/risk_jump/n54 , \t/a/condition/n1 , \t/a/risk_jump/n15 );  // PC.v(235)
  and \t/a/risk_jump/u32  (\t/a/risk_jump/n56 , \t/a/risk_jump/n54 , \t/memread_cs );  // PC.v(236)
  or \t/a/risk_jump/u33  (\t/a/risk_jump/n57 , \t/a/risk_jump/n24 , \t/a/risk_jump/n42 );  // PC.v(238)
  and \t/a/risk_jump/u34  (\t/a/risk_jump/n58 , \t/a/risk_jump/n56 , \t/a/risk_jump/n57 );  // PC.v(238)
  AL_MUX \t/a/risk_jump/u35  (
    .i0(\t/a/risk_jump/n58 ),
    .i1(1'b1),
    .sel(\t/a/risk_jump/n53 ),
    .o(\t/a/ID_jump_risk_block ));  // PC.v(240)
  and \t/a/risk_jump/u4  (\t/a/risk_jump/n5 , \t/a/condition/n1 , \t/a/n6 );  // PC.v(151)
  and \t/a/risk_jump/u5  (\t/a/risk_jump/MEM_risk , \t/a/risk_jump/n5 , \t/a/n7 );  // PC.v(152)
  and \t/a/risk_jump/u6  (\t/a/risk_jump/n8 , \t/a/condition/n1 , \t/a/n15 );  // PC.v(159)
  and \t/a/risk_jump/u7  (\t/a/risk_jump/WB_risk , \t/a/risk_jump/n8 , \t/a/n16 );  // PC.v(160)
  and \t/a/risk_jump/u8  (\t/a/risk_jump/n12 , \t/a/risk_jump/n10 , \t/a/risk_jump/n11 );  // PC.v(177)
  and \t/a/risk_jump/u9  (\t/a/risk_jump/n14 , \t/a/risk_jump/n12 , \t/a/risk_jump/n13 );  // PC.v(178)
  or \t/a/sel0_b10_sel  (\t/a/sel0_b10_sel_o , \t/a/n37 , \t/a/n36 );  // cpu.v(301)
  and \t/a/u10  (\t/a/n19 , \t/a/n17 , \t/a/n18 );  // cpu.v(245)
  and \t/a/u11  (\t/a/n21 , \t/a/n19 , \t/a/n20 );  // cpu.v(246)
  and \t/a/u12  (\t/a/n23 , \t/a/n21 , \t/a/n22 );  // cpu.v(247)
  and \t/a/u13  (\t/a/n25 , \t/a/n8 , \t/a/n24 );  // cpu.v(256)
  and \t/a/u14  (\t/a/n26 , \t/a/n25 , \t/a/n11 );  // cpu.v(257)
  and \t/a/u15  (\t/a/n27 , \t/a/n26 , \t/a/n13 );  // cpu.v(258)
  and \t/a/u17  (\t/a/n29 , \t/a/n19 , \t/a/n28 );  // cpu.v(263)
  and \t/a/u18  (\t/a/n31 , \t/a/n29 , \t/a/n30 );  // cpu.v(264)
  or \t/a/u19  (\t/a/n34 , \t/memread_cs , memwrite_cs);  // cpu.v(287)
  and \t/a/u2  (\t/a/n2 , \t/a/n0 , \t/a/n1 );  // cpu.v(179)
  or \t/a/u20  (\t/a/n33 , \t/a/n37 , \t/a/n32 );  // cpu.v(301)
  or \t/a/u21  (\t/a/n32 , \t/a/n36 , \t/a/n35 );  // cpu.v(301)
  or \t/a/u3  (\t/a/n5 , \t/a/n3 , \t/a/n4 );  // cpu.v(181)
  and \t/a/u4  (\t/a/ID_LW_block , \t/a/n2 , \t/a/n5 );  // cpu.v(181)
  and \t/a/u5  (\t/a/n8 , \t/a/n6 , \t/a/n7 );  // cpu.v(238)
  and \t/a/u6  (\t/a/n10 , \t/a/n8 , \t/a/n9 );  // cpu.v(239)
  and \t/a/u7  (\t/a/n12 , \t/a/n10 , \t/a/n11 );  // cpu.v(240)
  and \t/a/u8  (\t/a/n14 , \t/a/n12 , \t/a/n13 );  // cpu.v(241)
  and \t/a/u9  (\t/a/n17 , \t/a/n15 , \t/a/n16 );  // cpu.v(244)
  eq_w7 \t/a/unconditional/eq0  (
    .i0(\t/instruction [6:0]),
    .i1(7'b1101111),
    .o(\t/a/unconditional/n0 ));  // PC.v(100)
  eq_w7 \t/a/unconditional/eq1  (
    .i0(\t/instruction [6:0]),
    .i1(7'b0010111),
    .o(\t/a/unconditional/n1 ));  // PC.v(104)
  binary_mux_s1_w1 \t/a/unconditional/mux0_b20  (
    .i0(1'b0),
    .i1(\t/instruction [20]),
    .sel(\t/a/unconditional/n1 ),
    .o(\t/a/unconditional/n2 [20]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux0_b21  (
    .i0(1'b0),
    .i1(\t/instruction [21]),
    .sel(\t/a/unconditional/n1 ),
    .o(\t/a/unconditional/n2 [21]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux0_b22  (
    .i0(1'b0),
    .i1(\t/instruction [22]),
    .sel(\t/a/unconditional/n1 ),
    .o(\t/a/unconditional/n2 [22]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux0_b23  (
    .i0(1'b0),
    .i1(\t/instruction [23]),
    .sel(\t/a/unconditional/n1 ),
    .o(\t/a/unconditional/n2 [23]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux0_b24  (
    .i0(1'b0),
    .i1(\t/instruction [24]),
    .sel(\t/a/unconditional/n1 ),
    .o(\t/a/unconditional/n2 [24]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux0_b25  (
    .i0(1'b0),
    .i1(\t/instruction [25]),
    .sel(\t/a/unconditional/n1 ),
    .o(\t/a/unconditional/n2 [25]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux0_b26  (
    .i0(1'b0),
    .i1(\t/instruction [26]),
    .sel(\t/a/unconditional/n1 ),
    .o(\t/a/unconditional/n2 [26]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux0_b27  (
    .i0(1'b0),
    .i1(\t/instruction [27]),
    .sel(\t/a/unconditional/n1 ),
    .o(\t/a/unconditional/n2 [27]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux0_b28  (
    .i0(1'b0),
    .i1(\t/instruction [28]),
    .sel(\t/a/unconditional/n1 ),
    .o(\t/a/unconditional/n2 [28]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux0_b29  (
    .i0(1'b0),
    .i1(\t/instruction [29]),
    .sel(\t/a/unconditional/n1 ),
    .o(\t/a/unconditional/n2 [29]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux0_b30  (
    .i0(1'b0),
    .i1(\t/instruction [30]),
    .sel(\t/a/unconditional/n1 ),
    .o(\t/a/unconditional/n2 [30]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b1  (
    .i0(1'b0),
    .i1(\t/instruction [21]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [1]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b10  (
    .i0(1'b0),
    .i1(\t/instruction [30]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [10]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b11  (
    .i0(1'b0),
    .i1(\t/instruction [20]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [11]));  // PC.v(111)
  AL_MUX \t/a/unconditional/mux1_b12  (
    .i0(\t/instruction [12]),
    .i1(1'b0),
    .sel(\t/a/unconditional/mux1_b12_sel_is_0_o ),
    .o(\t/a/IF_skip_addr [12]));
  and \t/a/unconditional/mux1_b12_sel_is_0  (\t/a/unconditional/mux1_b12_sel_is_0_o , \t/a/unconditional/n0_neg , \t/a/unconditional/n1_neg );
  AL_MUX \t/a/unconditional/mux1_b13  (
    .i0(\t/instruction [13]),
    .i1(1'b0),
    .sel(\t/a/unconditional/mux1_b12_sel_is_0_o ),
    .o(\t/a/IF_skip_addr [13]));
  AL_MUX \t/a/unconditional/mux1_b14  (
    .i0(\t/instruction [14]),
    .i1(1'b0),
    .sel(\t/a/unconditional/mux1_b12_sel_is_0_o ),
    .o(\t/a/IF_skip_addr [14]));
  AL_MUX \t/a/unconditional/mux1_b15  (
    .i0(\t/instruction [15]),
    .i1(1'b0),
    .sel(\t/a/unconditional/mux1_b12_sel_is_0_o ),
    .o(\t/a/IF_skip_addr [15]));
  AL_MUX \t/a/unconditional/mux1_b16  (
    .i0(\t/instruction [16]),
    .i1(1'b0),
    .sel(\t/a/unconditional/mux1_b12_sel_is_0_o ),
    .o(\t/a/IF_skip_addr [16]));
  AL_MUX \t/a/unconditional/mux1_b17  (
    .i0(\t/instruction [17]),
    .i1(1'b0),
    .sel(\t/a/unconditional/mux1_b12_sel_is_0_o ),
    .o(\t/a/IF_skip_addr [17]));
  AL_MUX \t/a/unconditional/mux1_b18  (
    .i0(\t/instruction [18]),
    .i1(1'b0),
    .sel(\t/a/unconditional/mux1_b12_sel_is_0_o ),
    .o(\t/a/IF_skip_addr [18]));
  AL_MUX \t/a/unconditional/mux1_b19  (
    .i0(\t/instruction [19]),
    .i1(1'b0),
    .sel(\t/a/unconditional/mux1_b12_sel_is_0_o ),
    .o(\t/a/IF_skip_addr [19]));
  binary_mux_s1_w1 \t/a/unconditional/mux1_b2  (
    .i0(1'b0),
    .i1(\t/instruction [22]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [2]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b20  (
    .i0(\t/a/unconditional/n2 [20]),
    .i1(\t/instruction [31]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [20]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b21  (
    .i0(\t/a/unconditional/n2 [21]),
    .i1(\t/instruction [31]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [21]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b22  (
    .i0(\t/a/unconditional/n2 [22]),
    .i1(\t/instruction [31]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [22]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b23  (
    .i0(\t/a/unconditional/n2 [23]),
    .i1(\t/instruction [31]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [23]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b24  (
    .i0(\t/a/unconditional/n2 [24]),
    .i1(\t/instruction [31]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [24]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b25  (
    .i0(\t/a/unconditional/n2 [25]),
    .i1(\t/instruction [31]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [25]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b26  (
    .i0(\t/a/unconditional/n2 [26]),
    .i1(\t/instruction [31]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [26]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b27  (
    .i0(\t/a/unconditional/n2 [27]),
    .i1(\t/instruction [31]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [27]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b28  (
    .i0(\t/a/unconditional/n2 [28]),
    .i1(\t/instruction [31]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [28]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b29  (
    .i0(\t/a/unconditional/n2 [29]),
    .i1(\t/instruction [31]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [29]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b3  (
    .i0(1'b0),
    .i1(\t/instruction [23]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [3]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b30  (
    .i0(\t/a/unconditional/n2 [30]),
    .i1(\t/instruction [31]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [30]));  // PC.v(111)
  AL_MUX \t/a/unconditional/mux1_b31  (
    .i0(\t/instruction [31]),
    .i1(1'b0),
    .sel(\t/a/unconditional/mux1_b12_sel_is_0_o ),
    .o(\t/a/IF_skip_addr [31]));
  binary_mux_s1_w1 \t/a/unconditional/mux1_b4  (
    .i0(1'b0),
    .i1(\t/instruction [24]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [4]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b5  (
    .i0(1'b0),
    .i1(\t/instruction [25]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [5]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b6  (
    .i0(1'b0),
    .i1(\t/instruction [26]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [6]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b7  (
    .i0(1'b0),
    .i1(\t/instruction [27]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [7]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b8  (
    .i0(1'b0),
    .i1(\t/instruction [28]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [8]));  // PC.v(111)
  binary_mux_s1_w1 \t/a/unconditional/mux1_b9  (
    .i0(1'b0),
    .i1(\t/instruction [29]),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_addr [9]));  // PC.v(111)
  not \t/a/unconditional/n0_inv  (\t/a/unconditional/n0_neg , \t/a/unconditional/n0 );
  not \t/a/unconditional/n1_inv  (\t/a/unconditional/n1_neg , \t/a/unconditional/n1 );
  AL_MUX \t/a/unconditional/u2  (
    .i0(\t/a/unconditional/n1 ),
    .i1(1'b1),
    .sel(\t/a/unconditional/n0 ),
    .o(\t/a/IF_skip_cs ));  // PC.v(111)
  and \t/busarbitration/mux2_b0_sel_is_2  (\t/busarbitration/mux2_b0_sel_is_2_o , \t/a/instr/n1_neg , \t/a/mux3_b0_sel_is_1_o );
  and \t/busarbitration/mux2_b10_sel_is_2  (\t/busarbitration/mux2_b10_sel_is_2_o , \t/a/instr/n1_neg , \t/a/mux3_b10_sel_is_3_o );
  and \t/busarbitration/mux2_b16_sel_is_2  (\t/busarbitration/mux2_b16_sel_is_2_o , \t/a/instr/n1_neg , \t/a/mux3_b16_sel_is_3_o );
  binary_mux_s1_w1 \t/busarbitration/mux3_b0  (
    .i0(i_data[0]),
    .i1(\t/busarbitration/instruction [0]),
    .sel(\t/bus_block ),
    .o(\t/instruction [0]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b1  (
    .i0(i_data[1]),
    .i1(\t/busarbitration/instruction [1]),
    .sel(\t/bus_block ),
    .o(\t/instruction [1]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b10  (
    .i0(i_data[10]),
    .i1(\t/busarbitration/instruction [10]),
    .sel(\t/bus_block ),
    .o(\t/instruction [10]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b11  (
    .i0(i_data[11]),
    .i1(\t/busarbitration/instruction [11]),
    .sel(\t/bus_block ),
    .o(\t/instruction [11]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b12  (
    .i0(i_data[12]),
    .i1(\t/busarbitration/instruction [12]),
    .sel(\t/bus_block ),
    .o(\t/instruction [12]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b13  (
    .i0(i_data[13]),
    .i1(\t/busarbitration/instruction [13]),
    .sel(\t/bus_block ),
    .o(\t/instruction [13]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b14  (
    .i0(i_data[14]),
    .i1(\t/busarbitration/instruction [14]),
    .sel(\t/bus_block ),
    .o(\t/instruction [14]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b15  (
    .i0(i_data[15]),
    .i1(\t/busarbitration/instruction [15]),
    .sel(\t/bus_block ),
    .o(\t/instruction [15]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b16  (
    .i0(i_data[16]),
    .i1(\t/busarbitration/instruction [16]),
    .sel(\t/bus_block ),
    .o(\t/instruction [16]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b17  (
    .i0(i_data[17]),
    .i1(\t/busarbitration/instruction [17]),
    .sel(\t/bus_block ),
    .o(\t/instruction [17]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b18  (
    .i0(i_data[18]),
    .i1(\t/busarbitration/instruction [18]),
    .sel(\t/bus_block ),
    .o(\t/instruction [18]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b19  (
    .i0(i_data[19]),
    .i1(\t/busarbitration/instruction [19]),
    .sel(\t/bus_block ),
    .o(\t/instruction [19]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b2  (
    .i0(i_data[2]),
    .i1(\t/busarbitration/instruction [2]),
    .sel(\t/bus_block ),
    .o(\t/instruction [2]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b20  (
    .i0(i_data[20]),
    .i1(\t/busarbitration/instruction [20]),
    .sel(\t/bus_block ),
    .o(\t/instruction [20]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b21  (
    .i0(i_data[21]),
    .i1(\t/busarbitration/instruction [21]),
    .sel(\t/bus_block ),
    .o(\t/instruction [21]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b22  (
    .i0(i_data[22]),
    .i1(\t/busarbitration/instruction [22]),
    .sel(\t/bus_block ),
    .o(\t/instruction [22]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b23  (
    .i0(i_data[23]),
    .i1(\t/busarbitration/instruction [23]),
    .sel(\t/bus_block ),
    .o(\t/instruction [23]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b24  (
    .i0(i_data[24]),
    .i1(\t/busarbitration/instruction [24]),
    .sel(\t/bus_block ),
    .o(\t/instruction [24]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b25  (
    .i0(i_data[25]),
    .i1(\t/busarbitration/instruction [25]),
    .sel(\t/bus_block ),
    .o(\t/instruction [25]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b26  (
    .i0(i_data[26]),
    .i1(\t/busarbitration/instruction [26]),
    .sel(\t/bus_block ),
    .o(\t/instruction [26]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b27  (
    .i0(i_data[27]),
    .i1(\t/busarbitration/instruction [27]),
    .sel(\t/bus_block ),
    .o(\t/instruction [27]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b28  (
    .i0(i_data[28]),
    .i1(\t/busarbitration/instruction [28]),
    .sel(\t/bus_block ),
    .o(\t/instruction [28]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b29  (
    .i0(i_data[29]),
    .i1(\t/busarbitration/instruction [29]),
    .sel(\t/bus_block ),
    .o(\t/instruction [29]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b3  (
    .i0(i_data[3]),
    .i1(\t/busarbitration/instruction [3]),
    .sel(\t/bus_block ),
    .o(\t/instruction [3]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b30  (
    .i0(i_data[30]),
    .i1(\t/busarbitration/instruction [30]),
    .sel(\t/bus_block ),
    .o(\t/instruction [30]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b31  (
    .i0(i_data[31]),
    .i1(\t/busarbitration/instruction [31]),
    .sel(\t/bus_block ),
    .o(\t/instruction [31]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b4  (
    .i0(i_data[4]),
    .i1(\t/busarbitration/instruction [4]),
    .sel(\t/bus_block ),
    .o(\t/instruction [4]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b5  (
    .i0(i_data[5]),
    .i1(\t/busarbitration/instruction [5]),
    .sel(\t/bus_block ),
    .o(\t/instruction [5]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b6  (
    .i0(i_data[6]),
    .i1(\t/busarbitration/instruction [6]),
    .sel(\t/bus_block ),
    .o(\t/instruction [6]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b7  (
    .i0(i_data[7]),
    .i1(\t/busarbitration/instruction [7]),
    .sel(\t/bus_block ),
    .o(\t/instruction [7]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b8  (
    .i0(i_data[8]),
    .i1(\t/busarbitration/instruction [8]),
    .sel(\t/bus_block ),
    .o(\t/instruction [8]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux3_b9  (
    .i0(i_data[9]),
    .i1(\t/busarbitration/instruction [9]),
    .sel(\t/bus_block ),
    .o(\t/instruction [9]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b0  (
    .i0(\t/memstraddress [0]),
    .i1(\t/memaddress [0]),
    .sel(\t/bus_block ),
    .o(addr[0]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b1  (
    .i0(\t/memstraddress [1]),
    .i1(\t/memaddress [1]),
    .sel(\t/bus_block ),
    .o(addr[1]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b10  (
    .i0(\t/memstraddress [10]),
    .i1(\t/memaddress [10]),
    .sel(\t/bus_block ),
    .o(addr[10]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b11  (
    .i0(\t/memstraddress [11]),
    .i1(\t/memaddress [11]),
    .sel(\t/bus_block ),
    .o(addr[11]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b12  (
    .i0(\t/memstraddress [12]),
    .i1(\t/memaddress [12]),
    .sel(\t/bus_block ),
    .o(addr[12]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b13  (
    .i0(\t/memstraddress [13]),
    .i1(\t/memaddress [13]),
    .sel(\t/bus_block ),
    .o(addr[13]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b14  (
    .i0(\t/memstraddress [14]),
    .i1(\t/memaddress [14]),
    .sel(\t/bus_block ),
    .o(addr[14]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b15  (
    .i0(\t/memstraddress [15]),
    .i1(\t/memaddress [15]),
    .sel(\t/bus_block ),
    .o(addr[15]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b16  (
    .i0(\t/memstraddress [16]),
    .i1(\t/memaddress [16]),
    .sel(\t/bus_block ),
    .o(addr[16]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b17  (
    .i0(\t/memstraddress [17]),
    .i1(\t/memaddress [17]),
    .sel(\t/bus_block ),
    .o(addr[17]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b18  (
    .i0(\t/memstraddress [18]),
    .i1(\t/memaddress [18]),
    .sel(\t/bus_block ),
    .o(addr[18]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b19  (
    .i0(\t/memstraddress [19]),
    .i1(\t/memaddress [19]),
    .sel(\t/bus_block ),
    .o(addr[19]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b2  (
    .i0(\t/memstraddress [2]),
    .i1(\t/memaddress [2]),
    .sel(\t/bus_block ),
    .o(addr[2]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b20  (
    .i0(\t/memstraddress [20]),
    .i1(\t/memaddress [20]),
    .sel(\t/bus_block ),
    .o(addr[20]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b21  (
    .i0(\t/memstraddress [21]),
    .i1(\t/memaddress [21]),
    .sel(\t/bus_block ),
    .o(addr[21]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b22  (
    .i0(\t/memstraddress [22]),
    .i1(\t/memaddress [22]),
    .sel(\t/bus_block ),
    .o(addr[22]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b23  (
    .i0(\t/memstraddress [23]),
    .i1(\t/memaddress [23]),
    .sel(\t/bus_block ),
    .o(addr[23]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b24  (
    .i0(\t/memstraddress [24]),
    .i1(\t/memaddress [24]),
    .sel(\t/bus_block ),
    .o(addr[24]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b25  (
    .i0(\t/memstraddress [25]),
    .i1(\t/memaddress [25]),
    .sel(\t/bus_block ),
    .o(addr[25]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b26  (
    .i0(\t/memstraddress [26]),
    .i1(\t/memaddress [26]),
    .sel(\t/bus_block ),
    .o(addr[26]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b27  (
    .i0(\t/memstraddress [27]),
    .i1(\t/memaddress [27]),
    .sel(\t/bus_block ),
    .o(addr[27]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b28  (
    .i0(\t/memstraddress [28]),
    .i1(\t/memaddress [28]),
    .sel(\t/bus_block ),
    .o(addr[28]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b29  (
    .i0(\t/memstraddress [29]),
    .i1(\t/memaddress [29]),
    .sel(\t/bus_block ),
    .o(addr[29]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b3  (
    .i0(\t/memstraddress [3]),
    .i1(\t/memaddress [3]),
    .sel(\t/bus_block ),
    .o(addr[3]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b30  (
    .i0(\t/memstraddress [30]),
    .i1(\t/memaddress [30]),
    .sel(\t/bus_block ),
    .o(addr[30]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b31  (
    .i0(\t/memstraddress [31]),
    .i1(\t/memaddress [31]),
    .sel(\t/bus_block ),
    .o(addr[31]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b4  (
    .i0(\t/memstraddress [4]),
    .i1(\t/memaddress [4]),
    .sel(\t/bus_block ),
    .o(addr[4]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b5  (
    .i0(\t/memstraddress [5]),
    .i1(\t/memaddress [5]),
    .sel(\t/bus_block ),
    .o(addr[5]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b6  (
    .i0(\t/memstraddress [6]),
    .i1(\t/memaddress [6]),
    .sel(\t/bus_block ),
    .o(addr[6]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b7  (
    .i0(\t/memstraddress [7]),
    .i1(\t/memaddress [7]),
    .sel(\t/bus_block ),
    .o(addr[7]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b8  (
    .i0(\t/memstraddress [8]),
    .i1(\t/memaddress [8]),
    .sel(\t/bus_block ),
    .o(addr[8]));  // io.v(72)
  binary_mux_s1_w1 \t/busarbitration/mux4_b9  (
    .i0(\t/memstraddress [9]),
    .i1(\t/memaddress [9]),
    .sel(\t/bus_block ),
    .o(addr[9]));  // io.v(72)
  AL_MUX \t/busarbitration/mux5_b0  (
    .i0(1'b0),
    .i1(i_data[0]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [0]));
  and \t/busarbitration/mux5_b0_sel_is_3  (\t/busarbitration/mux5_b0_sel_is_3_o , \t/bus_block , \t/a/instr/n1 );
  AL_MUX \t/busarbitration/mux5_b1  (
    .i0(1'b0),
    .i1(i_data[1]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [1]));
  AL_MUX \t/busarbitration/mux5_b10  (
    .i0(1'b0),
    .i1(i_data[10]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [10]));
  AL_MUX \t/busarbitration/mux5_b11  (
    .i0(1'b0),
    .i1(i_data[11]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [11]));
  AL_MUX \t/busarbitration/mux5_b12  (
    .i0(1'b0),
    .i1(i_data[12]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [12]));
  AL_MUX \t/busarbitration/mux5_b13  (
    .i0(1'b0),
    .i1(i_data[13]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [13]));
  AL_MUX \t/busarbitration/mux5_b14  (
    .i0(1'b0),
    .i1(i_data[14]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [14]));
  AL_MUX \t/busarbitration/mux5_b15  (
    .i0(1'b0),
    .i1(i_data[15]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [15]));
  AL_MUX \t/busarbitration/mux5_b16  (
    .i0(1'b0),
    .i1(i_data[16]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [16]));
  AL_MUX \t/busarbitration/mux5_b17  (
    .i0(1'b0),
    .i1(i_data[17]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [17]));
  AL_MUX \t/busarbitration/mux5_b18  (
    .i0(1'b0),
    .i1(i_data[18]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [18]));
  AL_MUX \t/busarbitration/mux5_b19  (
    .i0(1'b0),
    .i1(i_data[19]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [19]));
  AL_MUX \t/busarbitration/mux5_b2  (
    .i0(1'b0),
    .i1(i_data[2]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [2]));
  AL_MUX \t/busarbitration/mux5_b20  (
    .i0(1'b0),
    .i1(i_data[20]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [20]));
  AL_MUX \t/busarbitration/mux5_b21  (
    .i0(1'b0),
    .i1(i_data[21]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [21]));
  AL_MUX \t/busarbitration/mux5_b22  (
    .i0(1'b0),
    .i1(i_data[22]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [22]));
  AL_MUX \t/busarbitration/mux5_b23  (
    .i0(1'b0),
    .i1(i_data[23]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [23]));
  AL_MUX \t/busarbitration/mux5_b24  (
    .i0(1'b0),
    .i1(i_data[24]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [24]));
  AL_MUX \t/busarbitration/mux5_b25  (
    .i0(1'b0),
    .i1(i_data[25]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [25]));
  AL_MUX \t/busarbitration/mux5_b26  (
    .i0(1'b0),
    .i1(i_data[26]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [26]));
  AL_MUX \t/busarbitration/mux5_b27  (
    .i0(1'b0),
    .i1(i_data[27]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [27]));
  AL_MUX \t/busarbitration/mux5_b28  (
    .i0(1'b0),
    .i1(i_data[28]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [28]));
  AL_MUX \t/busarbitration/mux5_b29  (
    .i0(1'b0),
    .i1(i_data[29]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [29]));
  AL_MUX \t/busarbitration/mux5_b3  (
    .i0(1'b0),
    .i1(i_data[3]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [3]));
  AL_MUX \t/busarbitration/mux5_b30  (
    .i0(1'b0),
    .i1(i_data[30]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [30]));
  AL_MUX \t/busarbitration/mux5_b31  (
    .i0(1'b0),
    .i1(i_data[31]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [31]));
  AL_MUX \t/busarbitration/mux5_b4  (
    .i0(1'b0),
    .i1(i_data[4]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [4]));
  AL_MUX \t/busarbitration/mux5_b5  (
    .i0(1'b0),
    .i1(i_data[5]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [5]));
  AL_MUX \t/busarbitration/mux5_b6  (
    .i0(1'b0),
    .i1(i_data[6]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [6]));
  AL_MUX \t/busarbitration/mux5_b7  (
    .i0(1'b0),
    .i1(i_data[7]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [7]));
  AL_MUX \t/busarbitration/mux5_b8  (
    .i0(1'b0),
    .i1(i_data[8]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [8]));
  AL_MUX \t/busarbitration/mux5_b9  (
    .i0(1'b0),
    .i1(i_data[9]),
    .sel(\t/busarbitration/mux5_b0_sel_is_3_o ),
    .o(\t/memreaddat [9]));
  AL_MUX \t/busarbitration/mux6_b0  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [0]),
    .sel(\t/busarbitration/mux6_b0_sel_is_3_o ),
    .o(o_data[0]));
  and \t/busarbitration/mux6_b0_sel_is_3  (\t/busarbitration/mux6_b0_sel_is_3_o , \t/bus_block , \t/busarbitration/mux2_b0_sel_is_2_o );
  AL_MUX \t/busarbitration/mux6_b1  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [1]),
    .sel(\t/busarbitration/mux6_b0_sel_is_3_o ),
    .o(o_data[1]));
  AL_MUX \t/busarbitration/mux6_b10  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [10]),
    .sel(\t/busarbitration/mux6_b10_sel_is_3_o ),
    .o(o_data[10]));
  and \t/busarbitration/mux6_b10_sel_is_3  (\t/busarbitration/mux6_b10_sel_is_3_o , \t/bus_block , \t/busarbitration/mux2_b10_sel_is_2_o );
  AL_MUX \t/busarbitration/mux6_b11  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [11]),
    .sel(\t/busarbitration/mux6_b10_sel_is_3_o ),
    .o(o_data[11]));
  AL_MUX \t/busarbitration/mux6_b12  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [12]),
    .sel(\t/busarbitration/mux6_b10_sel_is_3_o ),
    .o(o_data[12]));
  AL_MUX \t/busarbitration/mux6_b13  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [13]),
    .sel(\t/busarbitration/mux6_b10_sel_is_3_o ),
    .o(o_data[13]));
  AL_MUX \t/busarbitration/mux6_b14  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [14]),
    .sel(\t/busarbitration/mux6_b10_sel_is_3_o ),
    .o(o_data[14]));
  AL_MUX \t/busarbitration/mux6_b15  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [15]),
    .sel(\t/busarbitration/mux6_b10_sel_is_3_o ),
    .o(o_data[15]));
  AL_MUX \t/busarbitration/mux6_b16  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [16]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[16]));
  and \t/busarbitration/mux6_b16_sel_is_3  (\t/busarbitration/mux6_b16_sel_is_3_o , \t/bus_block , \t/busarbitration/mux2_b16_sel_is_2_o );
  AL_MUX \t/busarbitration/mux6_b17  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [17]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[17]));
  AL_MUX \t/busarbitration/mux6_b18  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [18]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[18]));
  AL_MUX \t/busarbitration/mux6_b19  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [19]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[19]));
  AL_MUX \t/busarbitration/mux6_b2  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [2]),
    .sel(\t/busarbitration/mux6_b0_sel_is_3_o ),
    .o(o_data[2]));
  AL_MUX \t/busarbitration/mux6_b20  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [20]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[20]));
  AL_MUX \t/busarbitration/mux6_b21  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [21]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[21]));
  AL_MUX \t/busarbitration/mux6_b22  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [22]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[22]));
  AL_MUX \t/busarbitration/mux6_b23  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [23]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[23]));
  AL_MUX \t/busarbitration/mux6_b24  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [24]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[24]));
  AL_MUX \t/busarbitration/mux6_b25  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [25]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[25]));
  AL_MUX \t/busarbitration/mux6_b26  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [26]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[26]));
  AL_MUX \t/busarbitration/mux6_b27  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [27]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[27]));
  AL_MUX \t/busarbitration/mux6_b28  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [28]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[28]));
  AL_MUX \t/busarbitration/mux6_b29  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [29]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[29]));
  AL_MUX \t/busarbitration/mux6_b3  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [3]),
    .sel(\t/busarbitration/mux6_b0_sel_is_3_o ),
    .o(o_data[3]));
  AL_MUX \t/busarbitration/mux6_b30  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [30]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[30]));
  AL_MUX \t/busarbitration/mux6_b31  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [31]),
    .sel(\t/busarbitration/mux6_b16_sel_is_3_o ),
    .o(o_data[31]));
  AL_MUX \t/busarbitration/mux6_b4  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [4]),
    .sel(\t/busarbitration/mux6_b0_sel_is_3_o ),
    .o(o_data[4]));
  AL_MUX \t/busarbitration/mux6_b5  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [5]),
    .sel(\t/busarbitration/mux6_b0_sel_is_3_o ),
    .o(o_data[5]));
  AL_MUX \t/busarbitration/mux6_b6  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [6]),
    .sel(\t/busarbitration/mux6_b0_sel_is_3_o ),
    .o(o_data[6]));
  AL_MUX \t/busarbitration/mux6_b7  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [7]),
    .sel(\t/busarbitration/mux6_b0_sel_is_3_o ),
    .o(o_data[7]));
  AL_MUX \t/busarbitration/mux6_b8  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [8]),
    .sel(\t/busarbitration/mux6_b10_sel_is_3_o ),
    .o(o_data[8]));
  AL_MUX \t/busarbitration/mux6_b9  (
    .i0(1'b0),
    .i1(\t/a/MEM_regdat2 [9]),
    .sel(\t/busarbitration/mux6_b10_sel_is_3_o ),
    .o(o_data[9]));
  ne_w1 \t/busarbitration/neq0  (
    .i0(\t/memread_cs ),
    .i1(1'b1),
    .o(\t/busarbitration/n1 ));  // io.v(45)
  ne_w1 \t/busarbitration/neq1  (
    .i0(memwrite_cs),
    .i1(1'b1),
    .o(\t/busarbitration/n2 ));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b0  (
    .clk(clock),
    .d(i_data[0]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [0]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b1  (
    .clk(clock),
    .d(i_data[1]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [1]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b10  (
    .clk(clock),
    .d(i_data[10]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [10]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b11  (
    .clk(clock),
    .d(i_data[11]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [11]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b12  (
    .clk(clock),
    .d(i_data[12]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [12]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b13  (
    .clk(clock),
    .d(i_data[13]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [13]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b14  (
    .clk(clock),
    .d(i_data[14]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [14]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b15  (
    .clk(clock),
    .d(i_data[15]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [15]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b16  (
    .clk(clock),
    .d(i_data[16]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [16]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b17  (
    .clk(clock),
    .d(i_data[17]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [17]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b18  (
    .clk(clock),
    .d(i_data[18]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [18]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b19  (
    .clk(clock),
    .d(i_data[19]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [19]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b2  (
    .clk(clock),
    .d(i_data[2]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [2]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b20  (
    .clk(clock),
    .d(i_data[20]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [20]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b21  (
    .clk(clock),
    .d(i_data[21]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [21]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b22  (
    .clk(clock),
    .d(i_data[22]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [22]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b23  (
    .clk(clock),
    .d(i_data[23]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [23]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b24  (
    .clk(clock),
    .d(i_data[24]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [24]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b25  (
    .clk(clock),
    .d(i_data[25]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [25]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b26  (
    .clk(clock),
    .d(i_data[26]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [26]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b27  (
    .clk(clock),
    .d(i_data[27]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [27]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b28  (
    .clk(clock),
    .d(i_data[28]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [28]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b29  (
    .clk(clock),
    .d(i_data[29]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [29]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b3  (
    .clk(clock),
    .d(i_data[3]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [3]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b30  (
    .clk(clock),
    .d(i_data[30]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [30]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b31  (
    .clk(clock),
    .d(i_data[31]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [31]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b4  (
    .clk(clock),
    .d(i_data[4]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [4]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b5  (
    .clk(clock),
    .d(i_data[5]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [5]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b6  (
    .clk(clock),
    .d(i_data[6]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [6]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b7  (
    .clk(clock),
    .d(i_data[7]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [7]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b8  (
    .clk(clock),
    .d(i_data[8]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [8]));  // io.v(45)
  reg_ar_as_w1 \t/busarbitration/reg0_b9  (
    .clk(clock),
    .d(i_data[9]),
    .en(\t/busarbitration/n3 ),
    .reset(~rst),
    .set(1'b0),
    .q(\t/busarbitration/instruction [9]));  // io.v(45)
  and \t/busarbitration/u4  (\t/busarbitration/n3 , \t/busarbitration/n1 , \t/busarbitration/n2 );  // io.v(45)
  or \t/busarbitration/u5  (\t/bus_block , \t/a/instr/n1 , n5);  // io.v(50)
  not \t/busarbitration/u6  (\t/instr_read , \t/bus_block );  // io.v(72)
  or \t/u0  (memread, \t/instr_read , \t/memread_cs );  // top2.v(21)
  and u2 (n1, memwrite_cs, n0);  // __top.v(51)
  and u4 (n7, n5, n6);  // __top.v(61)

endmodule 

module eq_w1
  (
  i0,
  i1,
  o
  );

  input i0;
  input i1;
  output o;

  wire xor_i0_i1_o;

  not none_diff (o, xor_i0_i1_o);
  xor xor_i0_i1 (xor_i0_i1_o, i0, i1);

endmodule 

module eq_w32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output o;

  wire or_or_or_or_or_xor_i_o;
  wire or_or_or_or_xor_i0$0_o;
  wire or_or_or_or_xor_i0$1_o;
  wire or_or_or_xor_i0$0$_i_o;
  wire or_or_or_xor_i0$16$__o;
  wire or_or_or_xor_i0$24$__o;
  wire or_or_or_xor_i0$8$_i_o;
  wire or_or_xor_i0$0$_i1$0_o;
  wire or_or_xor_i0$12$_i1$_o;
  wire or_or_xor_i0$16$_i1$_o;
  wire or_or_xor_i0$20$_i1$_o;
  wire or_or_xor_i0$24$_i1$_o;
  wire or_or_xor_i0$28$_i1$_o;
  wire or_or_xor_i0$4$_i1$4_o;
  wire or_or_xor_i0$8$_i1$8_o;
  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$10$_i1$10$_o;
  wire or_xor_i0$12$_i1$12$_o;
  wire or_xor_i0$14$_i1$14$_o;
  wire or_xor_i0$16$_i1$16$_o;
  wire or_xor_i0$18$_i1$18$_o;
  wire or_xor_i0$2$_i1$2$_o_o;
  wire or_xor_i0$20$_i1$20$_o;
  wire or_xor_i0$22$_i1$22$_o;
  wire or_xor_i0$24$_i1$24$_o;
  wire or_xor_i0$26$_i1$26$_o;
  wire or_xor_i0$28$_i1$28$_o;
  wire or_xor_i0$30$_i1$30$_o;
  wire or_xor_i0$4$_i1$4$_o_o;
  wire or_xor_i0$6$_i1$6$_o_o;
  wire or_xor_i0$8$_i1$8$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$10$_i1$10$_o;
  wire xor_i0$11$_i1$11$_o;
  wire xor_i0$12$_i1$12$_o;
  wire xor_i0$13$_i1$13$_o;
  wire xor_i0$14$_i1$14$_o;
  wire xor_i0$15$_i1$15$_o;
  wire xor_i0$16$_i1$16$_o;
  wire xor_i0$17$_i1$17$_o;
  wire xor_i0$18$_i1$18$_o;
  wire xor_i0$19$_i1$19$_o;
  wire xor_i0$2$_i1$2$_o;
  wire xor_i0$20$_i1$20$_o;
  wire xor_i0$21$_i1$21$_o;
  wire xor_i0$22$_i1$22$_o;
  wire xor_i0$23$_i1$23$_o;
  wire xor_i0$24$_i1$24$_o;
  wire xor_i0$25$_i1$25$_o;
  wire xor_i0$26$_i1$26$_o;
  wire xor_i0$27$_i1$27$_o;
  wire xor_i0$28$_i1$28$_o;
  wire xor_i0$29$_i1$29$_o;
  wire xor_i0$3$_i1$3$_o;
  wire xor_i0$30$_i1$30$_o;
  wire xor_i0$31$_i1$31$_o;
  wire xor_i0$4$_i1$4$_o;
  wire xor_i0$5$_i1$5$_o;
  wire xor_i0$6$_i1$6$_o;
  wire xor_i0$7$_i1$7$_o;
  wire xor_i0$8$_i1$8$_o;
  wire xor_i0$9$_i1$9$_o;

  not none_diff (o, or_or_or_or_or_xor_i_o);
  or or_or_or_or_or_xor_i (or_or_or_or_or_xor_i_o, or_or_or_or_xor_i0$0_o, or_or_or_or_xor_i0$1_o);
  or or_or_or_or_xor_i0$0 (or_or_or_or_xor_i0$0_o, or_or_or_xor_i0$0$_i_o, or_or_or_xor_i0$8$_i_o);
  or or_or_or_or_xor_i0$1 (or_or_or_or_xor_i0$1_o, or_or_or_xor_i0$16$__o, or_or_or_xor_i0$24$__o);
  or or_or_or_xor_i0$0$_i (or_or_or_xor_i0$0$_i_o, or_or_xor_i0$0$_i1$0_o, or_or_xor_i0$4$_i1$4_o);
  or or_or_or_xor_i0$16$_ (or_or_or_xor_i0$16$__o, or_or_xor_i0$16$_i1$_o, or_or_xor_i0$20$_i1$_o);
  or or_or_or_xor_i0$24$_ (or_or_or_xor_i0$24$__o, or_or_xor_i0$24$_i1$_o, or_or_xor_i0$28$_i1$_o);
  or or_or_or_xor_i0$8$_i (or_or_or_xor_i0$8$_i_o, or_or_xor_i0$8$_i1$8_o, or_or_xor_i0$12$_i1$_o);
  or or_or_xor_i0$0$_i1$0 (or_or_xor_i0$0$_i1$0_o, or_xor_i0$0$_i1$0$_o_o, or_xor_i0$2$_i1$2$_o_o);
  or or_or_xor_i0$12$_i1$ (or_or_xor_i0$12$_i1$_o, or_xor_i0$12$_i1$12$_o, or_xor_i0$14$_i1$14$_o);
  or or_or_xor_i0$16$_i1$ (or_or_xor_i0$16$_i1$_o, or_xor_i0$16$_i1$16$_o, or_xor_i0$18$_i1$18$_o);
  or or_or_xor_i0$20$_i1$ (or_or_xor_i0$20$_i1$_o, or_xor_i0$20$_i1$20$_o, or_xor_i0$22$_i1$22$_o);
  or or_or_xor_i0$24$_i1$ (or_or_xor_i0$24$_i1$_o, or_xor_i0$24$_i1$24$_o, or_xor_i0$26$_i1$26$_o);
  or or_or_xor_i0$28$_i1$ (or_or_xor_i0$28$_i1$_o, or_xor_i0$28$_i1$28$_o, or_xor_i0$30$_i1$30$_o);
  or or_or_xor_i0$4$_i1$4 (or_or_xor_i0$4$_i1$4_o, or_xor_i0$4$_i1$4$_o_o, or_xor_i0$6$_i1$6$_o_o);
  or or_or_xor_i0$8$_i1$8 (or_or_xor_i0$8$_i1$8_o, or_xor_i0$8$_i1$8$_o_o, or_xor_i0$10$_i1$10$_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, xor_i0$1$_i1$1$_o);
  or or_xor_i0$10$_i1$10$ (or_xor_i0$10$_i1$10$_o, xor_i0$10$_i1$10$_o, xor_i0$11$_i1$11$_o);
  or or_xor_i0$12$_i1$12$ (or_xor_i0$12$_i1$12$_o, xor_i0$12$_i1$12$_o, xor_i0$13$_i1$13$_o);
  or or_xor_i0$14$_i1$14$ (or_xor_i0$14$_i1$14$_o, xor_i0$14$_i1$14$_o, xor_i0$15$_i1$15$_o);
  or or_xor_i0$16$_i1$16$ (or_xor_i0$16$_i1$16$_o, xor_i0$16$_i1$16$_o, xor_i0$17$_i1$17$_o);
  or or_xor_i0$18$_i1$18$ (or_xor_i0$18$_i1$18$_o, xor_i0$18$_i1$18$_o, xor_i0$19$_i1$19$_o);
  or or_xor_i0$2$_i1$2$_o (or_xor_i0$2$_i1$2$_o_o, xor_i0$2$_i1$2$_o, xor_i0$3$_i1$3$_o);
  or or_xor_i0$20$_i1$20$ (or_xor_i0$20$_i1$20$_o, xor_i0$20$_i1$20$_o, xor_i0$21$_i1$21$_o);
  or or_xor_i0$22$_i1$22$ (or_xor_i0$22$_i1$22$_o, xor_i0$22$_i1$22$_o, xor_i0$23$_i1$23$_o);
  or or_xor_i0$24$_i1$24$ (or_xor_i0$24$_i1$24$_o, xor_i0$24$_i1$24$_o, xor_i0$25$_i1$25$_o);
  or or_xor_i0$26$_i1$26$ (or_xor_i0$26$_i1$26$_o, xor_i0$26$_i1$26$_o, xor_i0$27$_i1$27$_o);
  or or_xor_i0$28$_i1$28$ (or_xor_i0$28$_i1$28$_o, xor_i0$28$_i1$28$_o, xor_i0$29$_i1$29$_o);
  or or_xor_i0$30$_i1$30$ (or_xor_i0$30$_i1$30$_o, xor_i0$30$_i1$30$_o, xor_i0$31$_i1$31$_o);
  or or_xor_i0$4$_i1$4$_o (or_xor_i0$4$_i1$4$_o_o, xor_i0$4$_i1$4$_o, xor_i0$5$_i1$5$_o);
  or or_xor_i0$6$_i1$6$_o (or_xor_i0$6$_i1$6$_o_o, xor_i0$6$_i1$6$_o, xor_i0$7$_i1$7$_o);
  or or_xor_i0$8$_i1$8$_o (or_xor_i0$8$_i1$8$_o_o, xor_i0$8$_i1$8$_o, xor_i0$9$_i1$9$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (xor_i0$10$_i1$10$_o, i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (xor_i0$11$_i1$11$_o, i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (xor_i0$12$_i1$12$_o, i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (xor_i0$13$_i1$13$_o, i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (xor_i0$14$_i1$14$_o, i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (xor_i0$15$_i1$15$_o, i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (xor_i0$16$_i1$16$_o, i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (xor_i0$17$_i1$17$_o, i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (xor_i0$18$_i1$18$_o, i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (xor_i0$19$_i1$19$_o, i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (xor_i0$20$_i1$20$_o, i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (xor_i0$21$_i1$21$_o, i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (xor_i0$22$_i1$22$_o, i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (xor_i0$23$_i1$23$_o, i0[23], i1[23]);
  xor \xor_i0[24]_i1[24]  (xor_i0$24$_i1$24$_o, i0[24], i1[24]);
  xor \xor_i0[25]_i1[25]  (xor_i0$25$_i1$25$_o, i0[25], i1[25]);
  xor \xor_i0[26]_i1[26]  (xor_i0$26$_i1$26$_o, i0[26], i1[26]);
  xor \xor_i0[27]_i1[27]  (xor_i0$27$_i1$27$_o, i0[27], i1[27]);
  xor \xor_i0[28]_i1[28]  (xor_i0$28$_i1$28$_o, i0[28], i1[28]);
  xor \xor_i0[29]_i1[29]  (xor_i0$29$_i1$29$_o, i0[29], i1[29]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);
  xor \xor_i0[30]_i1[30]  (xor_i0$30$_i1$30$_o, i0[30], i1[30]);
  xor \xor_i0[31]_i1[31]  (xor_i0$31$_i1$31$_o, i0[31], i1[31]);
  xor \xor_i0[3]_i1[3]  (xor_i0$3$_i1$3$_o, i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (xor_i0$4$_i1$4$_o, i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (xor_i0$5$_i1$5$_o, i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (xor_i0$6$_i1$6$_o, i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (xor_i0$7$_i1$7$_o, i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (xor_i0$8$_i1$8$_o, i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (xor_i0$9$_i1$9$_o, i0[9], i1[9]);

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module lt_u32_u32
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [31:0] i0;
  input [31:0] i1;
  output o;

  wire [31:0] diff;
  wire diff_12_18;
  wire diff_19_26;
  wire diff_27_31;
  wire diff_6_11;
  wire less_12_18;
  wire \less_12_18_inst/diff_0 ;
  wire \less_12_18_inst/diff_1 ;
  wire \less_12_18_inst/diff_2 ;
  wire \less_12_18_inst/diff_3 ;
  wire \less_12_18_inst/diff_4 ;
  wire \less_12_18_inst/diff_5 ;
  wire \less_12_18_inst/diff_6 ;
  wire \less_12_18_inst/o_0 ;
  wire \less_12_18_inst/o_1 ;
  wire \less_12_18_inst/o_2 ;
  wire \less_12_18_inst/o_3 ;
  wire \less_12_18_inst/o_4 ;
  wire \less_12_18_inst/o_5 ;
  wire less_19_26;
  wire \less_19_26_inst/diff_0 ;
  wire \less_19_26_inst/diff_1 ;
  wire \less_19_26_inst/diff_2 ;
  wire \less_19_26_inst/diff_3 ;
  wire \less_19_26_inst/diff_4 ;
  wire \less_19_26_inst/diff_5 ;
  wire \less_19_26_inst/diff_6 ;
  wire \less_19_26_inst/diff_7 ;
  wire \less_19_26_inst/o_0 ;
  wire \less_19_26_inst/o_1 ;
  wire \less_19_26_inst/o_2 ;
  wire \less_19_26_inst/o_3 ;
  wire \less_19_26_inst/o_4 ;
  wire \less_19_26_inst/o_5 ;
  wire \less_19_26_inst/o_6 ;
  wire less_27_31;
  wire \less_27_31_inst/diff_0 ;
  wire \less_27_31_inst/diff_1 ;
  wire \less_27_31_inst/diff_2 ;
  wire \less_27_31_inst/diff_3 ;
  wire \less_27_31_inst/diff_4 ;
  wire \less_27_31_inst/o_0 ;
  wire \less_27_31_inst/o_1 ;
  wire \less_27_31_inst/o_2 ;
  wire \less_27_31_inst/o_3 ;
  wire less_6_11;
  wire \less_6_11_inst/diff_0 ;
  wire \less_6_11_inst/diff_1 ;
  wire \less_6_11_inst/diff_2 ;
  wire \less_6_11_inst/diff_3 ;
  wire \less_6_11_inst/diff_4 ;
  wire \less_6_11_inst/diff_5 ;
  wire \less_6_11_inst/o_0 ;
  wire \less_6_11_inst/o_1 ;
  wire \less_6_11_inst/o_2 ;
  wire \less_6_11_inst/o_3 ;
  wire \less_6_11_inst/o_4 ;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;
  wire o_6;
  wire o_7;
  wire o_8;

  or any_diff_12_18 (diff_12_18, diff[12], diff[13], diff[14], diff[15], diff[16], diff[17], diff[18]);
  or any_diff_19_26 (diff_19_26, diff[19], diff[20], diff[21], diff[22], diff[23], diff[24], diff[25], diff[26]);
  or any_diff_27_31 (diff_27_31, diff[27], diff[28], diff[29], diff[30], diff[31]);
  or any_diff_6_11 (diff_6_11, diff[6], diff[7], diff[8], diff[9], diff[10], diff[11]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_12 (diff[12], i0[12], i1[12]);
  xor diff_13 (diff[13], i0[13], i1[13]);
  xor diff_14 (diff[14], i0[14], i1[14]);
  xor diff_15 (diff[15], i0[15], i1[15]);
  xor diff_16 (diff[16], i0[16], i1[16]);
  xor diff_17 (diff[17], i0[17], i1[17]);
  xor diff_18 (diff[18], i0[18], i1[18]);
  xor diff_19 (diff[19], i0[19], i1[19]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_20 (diff[20], i0[20], i1[20]);
  xor diff_21 (diff[21], i0[21], i1[21]);
  xor diff_22 (diff[22], i0[22], i1[22]);
  xor diff_23 (diff[23], i0[23], i1[23]);
  xor diff_24 (diff[24], i0[24], i1[24]);
  xor diff_25 (diff[25], i0[25], i1[25]);
  xor diff_26 (diff[26], i0[26], i1[26]);
  xor diff_27 (diff[27], i0[27], i1[27]);
  xor diff_28 (diff[28], i0[28], i1[28]);
  xor diff_29 (diff[29], i0[29], i1[29]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_30 (diff[30], i0[30], i1[30]);
  xor diff_31 (diff[31], i0[31], i1[31]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_12_18_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[12]),
    .sel(\less_12_18_inst/diff_0 ),
    .o(\less_12_18_inst/o_0 ));
  AL_MUX \less_12_18_inst/mux_1  (
    .i0(\less_12_18_inst/o_0 ),
    .i1(i1[13]),
    .sel(\less_12_18_inst/diff_1 ),
    .o(\less_12_18_inst/o_1 ));
  AL_MUX \less_12_18_inst/mux_2  (
    .i0(\less_12_18_inst/o_1 ),
    .i1(i1[14]),
    .sel(\less_12_18_inst/diff_2 ),
    .o(\less_12_18_inst/o_2 ));
  AL_MUX \less_12_18_inst/mux_3  (
    .i0(\less_12_18_inst/o_2 ),
    .i1(i1[15]),
    .sel(\less_12_18_inst/diff_3 ),
    .o(\less_12_18_inst/o_3 ));
  AL_MUX \less_12_18_inst/mux_4  (
    .i0(\less_12_18_inst/o_3 ),
    .i1(i1[16]),
    .sel(\less_12_18_inst/diff_4 ),
    .o(\less_12_18_inst/o_4 ));
  AL_MUX \less_12_18_inst/mux_5  (
    .i0(\less_12_18_inst/o_4 ),
    .i1(i1[17]),
    .sel(\less_12_18_inst/diff_5 ),
    .o(\less_12_18_inst/o_5 ));
  AL_MUX \less_12_18_inst/mux_6  (
    .i0(\less_12_18_inst/o_5 ),
    .i1(i1[18]),
    .sel(\less_12_18_inst/diff_6 ),
    .o(less_12_18));
  xor \less_12_18_inst/xor_0  (\less_12_18_inst/diff_0 , i0[12], i1[12]);
  xor \less_12_18_inst/xor_1  (\less_12_18_inst/diff_1 , i0[13], i1[13]);
  xor \less_12_18_inst/xor_2  (\less_12_18_inst/diff_2 , i0[14], i1[14]);
  xor \less_12_18_inst/xor_3  (\less_12_18_inst/diff_3 , i0[15], i1[15]);
  xor \less_12_18_inst/xor_4  (\less_12_18_inst/diff_4 , i0[16], i1[16]);
  xor \less_12_18_inst/xor_5  (\less_12_18_inst/diff_5 , i0[17], i1[17]);
  xor \less_12_18_inst/xor_6  (\less_12_18_inst/diff_6 , i0[18], i1[18]);
  AL_MUX \less_19_26_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[19]),
    .sel(\less_19_26_inst/diff_0 ),
    .o(\less_19_26_inst/o_0 ));
  AL_MUX \less_19_26_inst/mux_1  (
    .i0(\less_19_26_inst/o_0 ),
    .i1(i1[20]),
    .sel(\less_19_26_inst/diff_1 ),
    .o(\less_19_26_inst/o_1 ));
  AL_MUX \less_19_26_inst/mux_2  (
    .i0(\less_19_26_inst/o_1 ),
    .i1(i1[21]),
    .sel(\less_19_26_inst/diff_2 ),
    .o(\less_19_26_inst/o_2 ));
  AL_MUX \less_19_26_inst/mux_3  (
    .i0(\less_19_26_inst/o_2 ),
    .i1(i1[22]),
    .sel(\less_19_26_inst/diff_3 ),
    .o(\less_19_26_inst/o_3 ));
  AL_MUX \less_19_26_inst/mux_4  (
    .i0(\less_19_26_inst/o_3 ),
    .i1(i1[23]),
    .sel(\less_19_26_inst/diff_4 ),
    .o(\less_19_26_inst/o_4 ));
  AL_MUX \less_19_26_inst/mux_5  (
    .i0(\less_19_26_inst/o_4 ),
    .i1(i1[24]),
    .sel(\less_19_26_inst/diff_5 ),
    .o(\less_19_26_inst/o_5 ));
  AL_MUX \less_19_26_inst/mux_6  (
    .i0(\less_19_26_inst/o_5 ),
    .i1(i1[25]),
    .sel(\less_19_26_inst/diff_6 ),
    .o(\less_19_26_inst/o_6 ));
  AL_MUX \less_19_26_inst/mux_7  (
    .i0(\less_19_26_inst/o_6 ),
    .i1(i1[26]),
    .sel(\less_19_26_inst/diff_7 ),
    .o(less_19_26));
  xor \less_19_26_inst/xor_0  (\less_19_26_inst/diff_0 , i0[19], i1[19]);
  xor \less_19_26_inst/xor_1  (\less_19_26_inst/diff_1 , i0[20], i1[20]);
  xor \less_19_26_inst/xor_2  (\less_19_26_inst/diff_2 , i0[21], i1[21]);
  xor \less_19_26_inst/xor_3  (\less_19_26_inst/diff_3 , i0[22], i1[22]);
  xor \less_19_26_inst/xor_4  (\less_19_26_inst/diff_4 , i0[23], i1[23]);
  xor \less_19_26_inst/xor_5  (\less_19_26_inst/diff_5 , i0[24], i1[24]);
  xor \less_19_26_inst/xor_6  (\less_19_26_inst/diff_6 , i0[25], i1[25]);
  xor \less_19_26_inst/xor_7  (\less_19_26_inst/diff_7 , i0[26], i1[26]);
  AL_MUX \less_27_31_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[27]),
    .sel(\less_27_31_inst/diff_0 ),
    .o(\less_27_31_inst/o_0 ));
  AL_MUX \less_27_31_inst/mux_1  (
    .i0(\less_27_31_inst/o_0 ),
    .i1(i1[28]),
    .sel(\less_27_31_inst/diff_1 ),
    .o(\less_27_31_inst/o_1 ));
  AL_MUX \less_27_31_inst/mux_2  (
    .i0(\less_27_31_inst/o_1 ),
    .i1(i1[29]),
    .sel(\less_27_31_inst/diff_2 ),
    .o(\less_27_31_inst/o_2 ));
  AL_MUX \less_27_31_inst/mux_3  (
    .i0(\less_27_31_inst/o_2 ),
    .i1(i1[30]),
    .sel(\less_27_31_inst/diff_3 ),
    .o(\less_27_31_inst/o_3 ));
  AL_MUX \less_27_31_inst/mux_4  (
    .i0(\less_27_31_inst/o_3 ),
    .i1(i1[31]),
    .sel(\less_27_31_inst/diff_4 ),
    .o(less_27_31));
  xor \less_27_31_inst/xor_0  (\less_27_31_inst/diff_0 , i0[27], i1[27]);
  xor \less_27_31_inst/xor_1  (\less_27_31_inst/diff_1 , i0[28], i1[28]);
  xor \less_27_31_inst/xor_2  (\less_27_31_inst/diff_2 , i0[29], i1[29]);
  xor \less_27_31_inst/xor_3  (\less_27_31_inst/diff_3 , i0[30], i1[30]);
  xor \less_27_31_inst/xor_4  (\less_27_31_inst/diff_4 , i0[31], i1[31]);
  AL_MUX \less_6_11_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_11_inst/diff_0 ),
    .o(\less_6_11_inst/o_0 ));
  AL_MUX \less_6_11_inst/mux_1  (
    .i0(\less_6_11_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_11_inst/diff_1 ),
    .o(\less_6_11_inst/o_1 ));
  AL_MUX \less_6_11_inst/mux_2  (
    .i0(\less_6_11_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_11_inst/diff_2 ),
    .o(\less_6_11_inst/o_2 ));
  AL_MUX \less_6_11_inst/mux_3  (
    .i0(\less_6_11_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_11_inst/diff_3 ),
    .o(\less_6_11_inst/o_3 ));
  AL_MUX \less_6_11_inst/mux_4  (
    .i0(\less_6_11_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_11_inst/diff_4 ),
    .o(\less_6_11_inst/o_4 ));
  AL_MUX \less_6_11_inst/mux_5  (
    .i0(\less_6_11_inst/o_4 ),
    .i1(i1[11]),
    .sel(\less_6_11_inst/diff_5 ),
    .o(less_6_11));
  xor \less_6_11_inst/xor_0  (\less_6_11_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_11_inst/xor_1  (\less_6_11_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_11_inst/xor_2  (\less_6_11_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_11_inst/xor_3  (\less_6_11_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_11_inst/xor_4  (\less_6_11_inst/diff_4 , i0[10], i1[10]);
  xor \less_6_11_inst/xor_5  (\less_6_11_inst/diff_5 , i0[11], i1[11]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_11),
    .sel(diff_6_11),
    .o(o_6));
  AL_MUX mux_7 (
    .i0(o_6),
    .i1(less_12_18),
    .sel(diff_12_18),
    .o(o_7));
  AL_MUX mux_8 (
    .i0(o_7),
    .i1(less_19_26),
    .sel(diff_19_26),
    .o(o_8));
  AL_MUX mux_9 (
    .i0(o_8),
    .i1(less_27_31),
    .sel(diff_27_31),
    .o(o));

endmodule 

module binary_mux_s1_w1
  (
  i0,
  i1,
  sel,
  o
  );

  input i0;
  input i1;
  input sel;
  output o;


  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel),
    .o(o));

endmodule 

module add_pu32_pu32_o32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [31:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module binary_mux_s4_w1
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  sel,
  o
  );

  input i0;
  input i1;
  input i10;
  input i11;
  input i12;
  input i13;
  input i14;
  input i15;
  input i2;
  input i3;
  input i4;
  input i5;
  input i6;
  input i7;
  input i8;
  input i9;
  input [3:0] sel;
  output o;

  wire  B0_0;
  wire  B0_1;
  wire  B0_2;
  wire  B0_3;
  wire  B0_4;
  wire  B0_5;
  wire  B0_6;
  wire  B0_7;
  wire  B1_0;
  wire  B1_1;
  wire  B1_2;
  wire  B1_3;
  wire  B2_0;
  wire  B2_1;

  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel[0]),
    .o(B0_0));
  AL_MUX al_mux_b0_0_1 (
    .i0(i2),
    .i1(i3),
    .sel(sel[0]),
    .o(B0_1));
  AL_MUX al_mux_b0_0_2 (
    .i0(i4),
    .i1(i5),
    .sel(sel[0]),
    .o(B0_2));
  AL_MUX al_mux_b0_0_3 (
    .i0(i6),
    .i1(i7),
    .sel(sel[0]),
    .o(B0_3));
  AL_MUX al_mux_b0_0_4 (
    .i0(i8),
    .i1(i9),
    .sel(sel[0]),
    .o(B0_4));
  AL_MUX al_mux_b0_0_5 (
    .i0(i10),
    .i1(i11),
    .sel(sel[0]),
    .o(B0_5));
  AL_MUX al_mux_b0_0_6 (
    .i0(i12),
    .i1(i13),
    .sel(sel[0]),
    .o(B0_6));
  AL_MUX al_mux_b0_0_7 (
    .i0(i14),
    .i1(i15),
    .sel(sel[0]),
    .o(B0_7));
  AL_MUX al_mux_b0_1_0 (
    .i0(B0_0),
    .i1(B0_1),
    .sel(sel[1]),
    .o(B1_0));
  AL_MUX al_mux_b0_1_1 (
    .i0(B0_2),
    .i1(B0_3),
    .sel(sel[1]),
    .o(B1_1));
  AL_MUX al_mux_b0_1_2 (
    .i0(B0_4),
    .i1(B0_5),
    .sel(sel[1]),
    .o(B1_2));
  AL_MUX al_mux_b0_1_3 (
    .i0(B0_6),
    .i1(B0_7),
    .sel(sel[1]),
    .o(B1_3));
  AL_MUX al_mux_b0_2_0 (
    .i0(B1_0),
    .i1(B1_1),
    .sel(sel[2]),
    .o(B2_0));
  AL_MUX al_mux_b0_2_1 (
    .i0(B1_2),
    .i1(B1_3),
    .sel(sel[2]),
    .o(B2_1));
  AL_MUX al_mux_b0_3_0 (
    .i0(B2_0),
    .i1(B2_1),
    .sel(sel[3]),
    .o(o));

endmodule 

module add_pu32_mu32_o32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [31:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb11;
  wire net_nb12;
  wire net_nb13;
  wire net_nb14;
  wire net_nb15;
  wire net_nb16;
  wire net_nb17;
  wire net_nb18;
  wire net_nb19;
  wire net_nb2;
  wire net_nb20;
  wire net_nb21;
  wire net_nb22;
  wire net_nb23;
  wire net_nb24;
  wire net_nb25;
  wire net_nb26;
  wire net_nb27;
  wire net_nb28;
  wire net_nb29;
  wire net_nb3;
  wire net_nb30;
  wire net_nb31;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_nb11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_nb12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_nb13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_nb14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_nb15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_nb16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_nb17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_nb18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_nb19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_nb20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_nb21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_nb22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_nb23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_nb24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_nb25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_nb26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_nb27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_nb28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_nb29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_nb30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_nb31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b11 (net_nb11, net_b11);
  not inv_b12 (net_nb12, net_b12);
  not inv_b13 (net_nb13, net_b13);
  not inv_b14 (net_nb14, net_b14);
  not inv_b15 (net_nb15, net_b15);
  not inv_b16 (net_nb16, net_b16);
  not inv_b17 (net_nb17, net_b17);
  not inv_b18 (net_nb18, net_b18);
  not inv_b19 (net_nb19, net_b19);
  not inv_b2 (net_nb2, net_b2);
  not inv_b20 (net_nb20, net_b20);
  not inv_b21 (net_nb21, net_b21);
  not inv_b22 (net_nb22, net_b22);
  not inv_b23 (net_nb23, net_b23);
  not inv_b24 (net_nb24, net_b24);
  not inv_b25 (net_nb25, net_b25);
  not inv_b26 (net_nb26, net_b26);
  not inv_b27 (net_nb27, net_b27);
  not inv_b28 (net_nb28, net_b28);
  not inv_b29 (net_nb29, net_b29);
  not inv_b3 (net_nb3, net_b3);
  not inv_b30 (net_nb30, net_b30);
  not inv_b31 (net_nb31, net_b31);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);

endmodule 

module eq_w7
  (
  i0,
  i1,
  o
  );

  input [6:0] i0;
  input [6:0] i1;
  output o;

  wire or_or_xor_i0$0$_i1$0_o;
  wire or_or_xor_i0$3$_i1$3_o;
  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$1$_i1$1$_o_o;
  wire or_xor_i0$3$_i1$3$_o_o;
  wire or_xor_i0$5$_i1$5$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$2$_i1$2$_o;
  wire xor_i0$3$_i1$3$_o;
  wire xor_i0$4$_i1$4$_o;
  wire xor_i0$5$_i1$5$_o;
  wire xor_i0$6$_i1$6$_o;

  not none_diff (o, or_or_xor_i0$0$_i1$0_o);
  or or_or_xor_i0$0$_i1$0 (or_or_xor_i0$0$_i1$0_o, or_xor_i0$0$_i1$0$_o_o, or_or_xor_i0$3$_i1$3_o);
  or or_or_xor_i0$3$_i1$3 (or_or_xor_i0$3$_i1$3_o, or_xor_i0$3$_i1$3$_o_o, or_xor_i0$5$_i1$5$_o_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, or_xor_i0$1$_i1$1$_o_o);
  or or_xor_i0$1$_i1$1$_o (or_xor_i0$1$_i1$1$_o_o, xor_i0$1$_i1$1$_o, xor_i0$2$_i1$2$_o);
  or or_xor_i0$3$_i1$3$_o (or_xor_i0$3$_i1$3$_o_o, xor_i0$3$_i1$3$_o, xor_i0$4$_i1$4$_o);
  or or_xor_i0$5$_i1$5$_o (or_xor_i0$5$_i1$5$_o_o, xor_i0$5$_i1$5$_o, xor_i0$6$_i1$6$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (xor_i0$3$_i1$3$_o, i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (xor_i0$4$_i1$4$_o, i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (xor_i0$5$_i1$5$_o, i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (xor_i0$6$_i1$6$_o, i0[6], i1[6]);

endmodule 

module eq_w3
  (
  i0,
  i1,
  o
  );

  input [2:0] i0;
  input [2:0] i1;
  output o;

  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$1$_i1$1$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$2$_i1$2$_o;

  not none_diff (o, or_xor_i0$0$_i1$0$_o_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, or_xor_i0$1$_i1$1$_o_o);
  or or_xor_i0$1$_i1$1$_o (or_xor_i0$1$_i1$1$_o_o, xor_i0$1$_i1$1$_o, xor_i0$2$_i1$2$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);

endmodule 

module binary_mux_s2_w1
  (
  i0,
  i1,
  i2,
  i3,
  sel,
  o
  );

  input i0;
  input i1;
  input i2;
  input i3;
  input [1:0] sel;
  output o;

  wire  B0_0;
  wire  B0_1;

  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel[0]),
    .o(B0_0));
  AL_MUX al_mux_b0_0_1 (
    .i0(i2),
    .i1(i3),
    .sel(sel[0]),
    .o(B0_1));
  AL_MUX al_mux_b0_1_0 (
    .i0(B0_0),
    .i1(B0_1),
    .sel(sel[1]),
    .o(o));

endmodule 

module lt_u31_u31
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [30:0] i0;
  input [30:0] i1;
  output o;

  wire [30:0] diff;
  wire diff_12_18;
  wire diff_19_26;
  wire diff_27_30;
  wire diff_6_11;
  wire less_12_18;
  wire \less_12_18_inst/diff_0 ;
  wire \less_12_18_inst/diff_1 ;
  wire \less_12_18_inst/diff_2 ;
  wire \less_12_18_inst/diff_3 ;
  wire \less_12_18_inst/diff_4 ;
  wire \less_12_18_inst/diff_5 ;
  wire \less_12_18_inst/diff_6 ;
  wire \less_12_18_inst/o_0 ;
  wire \less_12_18_inst/o_1 ;
  wire \less_12_18_inst/o_2 ;
  wire \less_12_18_inst/o_3 ;
  wire \less_12_18_inst/o_4 ;
  wire \less_12_18_inst/o_5 ;
  wire less_19_26;
  wire \less_19_26_inst/diff_0 ;
  wire \less_19_26_inst/diff_1 ;
  wire \less_19_26_inst/diff_2 ;
  wire \less_19_26_inst/diff_3 ;
  wire \less_19_26_inst/diff_4 ;
  wire \less_19_26_inst/diff_5 ;
  wire \less_19_26_inst/diff_6 ;
  wire \less_19_26_inst/diff_7 ;
  wire \less_19_26_inst/o_0 ;
  wire \less_19_26_inst/o_1 ;
  wire \less_19_26_inst/o_2 ;
  wire \less_19_26_inst/o_3 ;
  wire \less_19_26_inst/o_4 ;
  wire \less_19_26_inst/o_5 ;
  wire \less_19_26_inst/o_6 ;
  wire less_27_30;
  wire \less_27_30_inst/diff_0 ;
  wire \less_27_30_inst/diff_1 ;
  wire \less_27_30_inst/diff_2 ;
  wire \less_27_30_inst/diff_3 ;
  wire \less_27_30_inst/o_0 ;
  wire \less_27_30_inst/o_1 ;
  wire \less_27_30_inst/o_2 ;
  wire less_6_11;
  wire \less_6_11_inst/diff_0 ;
  wire \less_6_11_inst/diff_1 ;
  wire \less_6_11_inst/diff_2 ;
  wire \less_6_11_inst/diff_3 ;
  wire \less_6_11_inst/diff_4 ;
  wire \less_6_11_inst/diff_5 ;
  wire \less_6_11_inst/o_0 ;
  wire \less_6_11_inst/o_1 ;
  wire \less_6_11_inst/o_2 ;
  wire \less_6_11_inst/o_3 ;
  wire \less_6_11_inst/o_4 ;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;
  wire o_6;
  wire o_7;
  wire o_8;

  or any_diff_12_18 (diff_12_18, diff[12], diff[13], diff[14], diff[15], diff[16], diff[17], diff[18]);
  or any_diff_19_26 (diff_19_26, diff[19], diff[20], diff[21], diff[22], diff[23], diff[24], diff[25], diff[26]);
  or any_diff_27_30 (diff_27_30, diff[27], diff[28], diff[29], diff[30]);
  or any_diff_6_11 (diff_6_11, diff[6], diff[7], diff[8], diff[9], diff[10], diff[11]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_12 (diff[12], i0[12], i1[12]);
  xor diff_13 (diff[13], i0[13], i1[13]);
  xor diff_14 (diff[14], i0[14], i1[14]);
  xor diff_15 (diff[15], i0[15], i1[15]);
  xor diff_16 (diff[16], i0[16], i1[16]);
  xor diff_17 (diff[17], i0[17], i1[17]);
  xor diff_18 (diff[18], i0[18], i1[18]);
  xor diff_19 (diff[19], i0[19], i1[19]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_20 (diff[20], i0[20], i1[20]);
  xor diff_21 (diff[21], i0[21], i1[21]);
  xor diff_22 (diff[22], i0[22], i1[22]);
  xor diff_23 (diff[23], i0[23], i1[23]);
  xor diff_24 (diff[24], i0[24], i1[24]);
  xor diff_25 (diff[25], i0[25], i1[25]);
  xor diff_26 (diff[26], i0[26], i1[26]);
  xor diff_27 (diff[27], i0[27], i1[27]);
  xor diff_28 (diff[28], i0[28], i1[28]);
  xor diff_29 (diff[29], i0[29], i1[29]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_30 (diff[30], i0[30], i1[30]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_12_18_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[12]),
    .sel(\less_12_18_inst/diff_0 ),
    .o(\less_12_18_inst/o_0 ));
  AL_MUX \less_12_18_inst/mux_1  (
    .i0(\less_12_18_inst/o_0 ),
    .i1(i1[13]),
    .sel(\less_12_18_inst/diff_1 ),
    .o(\less_12_18_inst/o_1 ));
  AL_MUX \less_12_18_inst/mux_2  (
    .i0(\less_12_18_inst/o_1 ),
    .i1(i1[14]),
    .sel(\less_12_18_inst/diff_2 ),
    .o(\less_12_18_inst/o_2 ));
  AL_MUX \less_12_18_inst/mux_3  (
    .i0(\less_12_18_inst/o_2 ),
    .i1(i1[15]),
    .sel(\less_12_18_inst/diff_3 ),
    .o(\less_12_18_inst/o_3 ));
  AL_MUX \less_12_18_inst/mux_4  (
    .i0(\less_12_18_inst/o_3 ),
    .i1(i1[16]),
    .sel(\less_12_18_inst/diff_4 ),
    .o(\less_12_18_inst/o_4 ));
  AL_MUX \less_12_18_inst/mux_5  (
    .i0(\less_12_18_inst/o_4 ),
    .i1(i1[17]),
    .sel(\less_12_18_inst/diff_5 ),
    .o(\less_12_18_inst/o_5 ));
  AL_MUX \less_12_18_inst/mux_6  (
    .i0(\less_12_18_inst/o_5 ),
    .i1(i1[18]),
    .sel(\less_12_18_inst/diff_6 ),
    .o(less_12_18));
  xor \less_12_18_inst/xor_0  (\less_12_18_inst/diff_0 , i0[12], i1[12]);
  xor \less_12_18_inst/xor_1  (\less_12_18_inst/diff_1 , i0[13], i1[13]);
  xor \less_12_18_inst/xor_2  (\less_12_18_inst/diff_2 , i0[14], i1[14]);
  xor \less_12_18_inst/xor_3  (\less_12_18_inst/diff_3 , i0[15], i1[15]);
  xor \less_12_18_inst/xor_4  (\less_12_18_inst/diff_4 , i0[16], i1[16]);
  xor \less_12_18_inst/xor_5  (\less_12_18_inst/diff_5 , i0[17], i1[17]);
  xor \less_12_18_inst/xor_6  (\less_12_18_inst/diff_6 , i0[18], i1[18]);
  AL_MUX \less_19_26_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[19]),
    .sel(\less_19_26_inst/diff_0 ),
    .o(\less_19_26_inst/o_0 ));
  AL_MUX \less_19_26_inst/mux_1  (
    .i0(\less_19_26_inst/o_0 ),
    .i1(i1[20]),
    .sel(\less_19_26_inst/diff_1 ),
    .o(\less_19_26_inst/o_1 ));
  AL_MUX \less_19_26_inst/mux_2  (
    .i0(\less_19_26_inst/o_1 ),
    .i1(i1[21]),
    .sel(\less_19_26_inst/diff_2 ),
    .o(\less_19_26_inst/o_2 ));
  AL_MUX \less_19_26_inst/mux_3  (
    .i0(\less_19_26_inst/o_2 ),
    .i1(i1[22]),
    .sel(\less_19_26_inst/diff_3 ),
    .o(\less_19_26_inst/o_3 ));
  AL_MUX \less_19_26_inst/mux_4  (
    .i0(\less_19_26_inst/o_3 ),
    .i1(i1[23]),
    .sel(\less_19_26_inst/diff_4 ),
    .o(\less_19_26_inst/o_4 ));
  AL_MUX \less_19_26_inst/mux_5  (
    .i0(\less_19_26_inst/o_4 ),
    .i1(i1[24]),
    .sel(\less_19_26_inst/diff_5 ),
    .o(\less_19_26_inst/o_5 ));
  AL_MUX \less_19_26_inst/mux_6  (
    .i0(\less_19_26_inst/o_5 ),
    .i1(i1[25]),
    .sel(\less_19_26_inst/diff_6 ),
    .o(\less_19_26_inst/o_6 ));
  AL_MUX \less_19_26_inst/mux_7  (
    .i0(\less_19_26_inst/o_6 ),
    .i1(i1[26]),
    .sel(\less_19_26_inst/diff_7 ),
    .o(less_19_26));
  xor \less_19_26_inst/xor_0  (\less_19_26_inst/diff_0 , i0[19], i1[19]);
  xor \less_19_26_inst/xor_1  (\less_19_26_inst/diff_1 , i0[20], i1[20]);
  xor \less_19_26_inst/xor_2  (\less_19_26_inst/diff_2 , i0[21], i1[21]);
  xor \less_19_26_inst/xor_3  (\less_19_26_inst/diff_3 , i0[22], i1[22]);
  xor \less_19_26_inst/xor_4  (\less_19_26_inst/diff_4 , i0[23], i1[23]);
  xor \less_19_26_inst/xor_5  (\less_19_26_inst/diff_5 , i0[24], i1[24]);
  xor \less_19_26_inst/xor_6  (\less_19_26_inst/diff_6 , i0[25], i1[25]);
  xor \less_19_26_inst/xor_7  (\less_19_26_inst/diff_7 , i0[26], i1[26]);
  AL_MUX \less_27_30_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[27]),
    .sel(\less_27_30_inst/diff_0 ),
    .o(\less_27_30_inst/o_0 ));
  AL_MUX \less_27_30_inst/mux_1  (
    .i0(\less_27_30_inst/o_0 ),
    .i1(i1[28]),
    .sel(\less_27_30_inst/diff_1 ),
    .o(\less_27_30_inst/o_1 ));
  AL_MUX \less_27_30_inst/mux_2  (
    .i0(\less_27_30_inst/o_1 ),
    .i1(i1[29]),
    .sel(\less_27_30_inst/diff_2 ),
    .o(\less_27_30_inst/o_2 ));
  AL_MUX \less_27_30_inst/mux_3  (
    .i0(\less_27_30_inst/o_2 ),
    .i1(i1[30]),
    .sel(\less_27_30_inst/diff_3 ),
    .o(less_27_30));
  xor \less_27_30_inst/xor_0  (\less_27_30_inst/diff_0 , i0[27], i1[27]);
  xor \less_27_30_inst/xor_1  (\less_27_30_inst/diff_1 , i0[28], i1[28]);
  xor \less_27_30_inst/xor_2  (\less_27_30_inst/diff_2 , i0[29], i1[29]);
  xor \less_27_30_inst/xor_3  (\less_27_30_inst/diff_3 , i0[30], i1[30]);
  AL_MUX \less_6_11_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_11_inst/diff_0 ),
    .o(\less_6_11_inst/o_0 ));
  AL_MUX \less_6_11_inst/mux_1  (
    .i0(\less_6_11_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_11_inst/diff_1 ),
    .o(\less_6_11_inst/o_1 ));
  AL_MUX \less_6_11_inst/mux_2  (
    .i0(\less_6_11_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_11_inst/diff_2 ),
    .o(\less_6_11_inst/o_2 ));
  AL_MUX \less_6_11_inst/mux_3  (
    .i0(\less_6_11_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_11_inst/diff_3 ),
    .o(\less_6_11_inst/o_3 ));
  AL_MUX \less_6_11_inst/mux_4  (
    .i0(\less_6_11_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_11_inst/diff_4 ),
    .o(\less_6_11_inst/o_4 ));
  AL_MUX \less_6_11_inst/mux_5  (
    .i0(\less_6_11_inst/o_4 ),
    .i1(i1[11]),
    .sel(\less_6_11_inst/diff_5 ),
    .o(less_6_11));
  xor \less_6_11_inst/xor_0  (\less_6_11_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_11_inst/xor_1  (\less_6_11_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_11_inst/xor_2  (\less_6_11_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_11_inst/xor_3  (\less_6_11_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_11_inst/xor_4  (\less_6_11_inst/diff_4 , i0[10], i1[10]);
  xor \less_6_11_inst/xor_5  (\less_6_11_inst/diff_5 , i0[11], i1[11]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_11),
    .sel(diff_6_11),
    .o(o_6));
  AL_MUX mux_7 (
    .i0(o_6),
    .i1(less_12_18),
    .sel(diff_12_18),
    .o(o_7));
  AL_MUX mux_8 (
    .i0(o_7),
    .i1(less_19_26),
    .sel(diff_19_26),
    .o(o_8));
  AL_MUX mux_9 (
    .i0(o_8),
    .i1(less_27_30),
    .sel(diff_27_30),
    .o(o));

endmodule 

module binary_mux_s3_w1
  (
  i0,
  i1,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  sel,
  o
  );

  input i0;
  input i1;
  input i2;
  input i3;
  input i4;
  input i5;
  input i6;
  input i7;
  input [2:0] sel;
  output o;

  wire  B0_0;
  wire  B0_1;
  wire  B0_2;
  wire  B0_3;
  wire  B1_0;
  wire  B1_1;

  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel[0]),
    .o(B0_0));
  AL_MUX al_mux_b0_0_1 (
    .i0(i2),
    .i1(i3),
    .sel(sel[0]),
    .o(B0_1));
  AL_MUX al_mux_b0_0_2 (
    .i0(i4),
    .i1(i5),
    .sel(sel[0]),
    .o(B0_2));
  AL_MUX al_mux_b0_0_3 (
    .i0(i6),
    .i1(i7),
    .sel(sel[0]),
    .o(B0_3));
  AL_MUX al_mux_b0_1_0 (
    .i0(B0_0),
    .i1(B0_1),
    .sel(sel[1]),
    .o(B1_0));
  AL_MUX al_mux_b0_1_1 (
    .i0(B0_2),
    .i1(B0_3),
    .sel(sel[1]),
    .o(B1_1));
  AL_MUX al_mux_b0_2_0 (
    .i0(B1_0),
    .i1(B1_1),
    .sel(sel[2]),
    .o(o));

endmodule 

module ne_w32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output o;

  wire [31:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3], diff[4], diff[5], diff[6], diff[7], diff[8], diff[9], diff[10], diff[11], diff[12], diff[13], diff[14], diff[15], diff[16], diff[17], diff[18], diff[19], diff[20], diff[21], diff[22], diff[23], diff[24], diff[25], diff[26], diff[27], diff[28], diff[29], diff[30], diff[31]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_12 (diff[12], i0[12], i1[12]);
  xor diff_13 (diff[13], i0[13], i1[13]);
  xor diff_14 (diff[14], i0[14], i1[14]);
  xor diff_15 (diff[15], i0[15], i1[15]);
  xor diff_16 (diff[16], i0[16], i1[16]);
  xor diff_17 (diff[17], i0[17], i1[17]);
  xor diff_18 (diff[18], i0[18], i1[18]);
  xor diff_19 (diff[19], i0[19], i1[19]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_20 (diff[20], i0[20], i1[20]);
  xor diff_21 (diff[21], i0[21], i1[21]);
  xor diff_22 (diff[22], i0[22], i1[22]);
  xor diff_23 (diff[23], i0[23], i1[23]);
  xor diff_24 (diff[24], i0[24], i1[24]);
  xor diff_25 (diff[25], i0[25], i1[25]);
  xor diff_26 (diff[26], i0[26], i1[26]);
  xor diff_27 (diff[27], i0[27], i1[27]);
  xor diff_28 (diff[28], i0[28], i1[28]);
  xor diff_29 (diff[29], i0[29], i1[29]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_30 (diff[30], i0[30], i1[30]);
  xor diff_31 (diff[31], i0[31], i1[31]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);

endmodule 

module eq_w5
  (
  i0,
  i1,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  output o;

  wire or_or_xor_i0$0$_i1$0_o;
  wire or_xor_i0$0$_i1$0$_o_o;
  wire or_xor_i0$2$_i1$2$_o_o;
  wire or_xor_i0$3$_i1$3$_o_o;
  wire xor_i0$0$_i1$0$_o;
  wire xor_i0$1$_i1$1$_o;
  wire xor_i0$2$_i1$2$_o;
  wire xor_i0$3$_i1$3$_o;
  wire xor_i0$4$_i1$4$_o;

  not none_diff (o, or_or_xor_i0$0$_i1$0_o);
  or or_or_xor_i0$0$_i1$0 (or_or_xor_i0$0$_i1$0_o, or_xor_i0$0$_i1$0$_o_o, or_xor_i0$2$_i1$2$_o_o);
  or or_xor_i0$0$_i1$0$_o (or_xor_i0$0$_i1$0$_o_o, xor_i0$0$_i1$0$_o, xor_i0$1$_i1$1$_o);
  or or_xor_i0$2$_i1$2$_o (or_xor_i0$2$_i1$2$_o_o, xor_i0$2$_i1$2$_o, or_xor_i0$3$_i1$3$_o_o);
  or or_xor_i0$3$_i1$3$_o (or_xor_i0$3$_i1$3$_o_o, xor_i0$3$_i1$3$_o, xor_i0$4$_i1$4$_o);
  xor \xor_i0[0]_i1[0]  (xor_i0$0$_i1$0$_o, i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (xor_i0$1$_i1$1$_o, i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (xor_i0$2$_i1$2$_o, i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (xor_i0$3$_i1$3$_o, i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (xor_i0$4$_i1$4$_o, i0[4], i1[4]);

endmodule 

module add_pu30_pu30_o30
  (
  i0,
  i1,
  o
  );

  input [29:0] i0;
  input [29:0] i1;
  output [29:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module ne_w7
  (
  i0,
  i1,
  o
  );

  input [6:0] i0;
  input [6:0] i1;
  output o;

  wire [6:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3], diff[4], diff[5], diff[6]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);

endmodule 

module ne_w5
  (
  i0,
  i1,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  output o;

  wire [4:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3], diff[4]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);

endmodule 

module binary_mux_s5_w1
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i16,
  i17,
  i18,
  i19,
  i2,
  i20,
  i21,
  i22,
  i23,
  i24,
  i25,
  i26,
  i27,
  i28,
  i29,
  i3,
  i30,
  i31,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  sel,
  o
  );

  input i0;
  input i1;
  input i10;
  input i11;
  input i12;
  input i13;
  input i14;
  input i15;
  input i16;
  input i17;
  input i18;
  input i19;
  input i2;
  input i20;
  input i21;
  input i22;
  input i23;
  input i24;
  input i25;
  input i26;
  input i27;
  input i28;
  input i29;
  input i3;
  input i30;
  input i31;
  input i4;
  input i5;
  input i6;
  input i7;
  input i8;
  input i9;
  input [4:0] sel;
  output o;

  wire  B0_0;
  wire  B0_1;
  wire  B0_10;
  wire  B0_11;
  wire  B0_12;
  wire  B0_13;
  wire  B0_14;
  wire  B0_15;
  wire  B0_2;
  wire  B0_3;
  wire  B0_4;
  wire  B0_5;
  wire  B0_6;
  wire  B0_7;
  wire  B0_8;
  wire  B0_9;
  wire  B1_0;
  wire  B1_1;
  wire  B1_2;
  wire  B1_3;
  wire  B1_4;
  wire  B1_5;
  wire  B1_6;
  wire  B1_7;
  wire  B2_0;
  wire  B2_1;
  wire  B2_2;
  wire  B2_3;
  wire  B3_0;
  wire  B3_1;

  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel[0]),
    .o(B0_0));
  AL_MUX al_mux_b0_0_1 (
    .i0(i2),
    .i1(i3),
    .sel(sel[0]),
    .o(B0_1));
  AL_MUX al_mux_b0_0_10 (
    .i0(i20),
    .i1(i21),
    .sel(sel[0]),
    .o(B0_10));
  AL_MUX al_mux_b0_0_11 (
    .i0(i22),
    .i1(i23),
    .sel(sel[0]),
    .o(B0_11));
  AL_MUX al_mux_b0_0_12 (
    .i0(i24),
    .i1(i25),
    .sel(sel[0]),
    .o(B0_12));
  AL_MUX al_mux_b0_0_13 (
    .i0(i26),
    .i1(i27),
    .sel(sel[0]),
    .o(B0_13));
  AL_MUX al_mux_b0_0_14 (
    .i0(i28),
    .i1(i29),
    .sel(sel[0]),
    .o(B0_14));
  AL_MUX al_mux_b0_0_15 (
    .i0(i30),
    .i1(i31),
    .sel(sel[0]),
    .o(B0_15));
  AL_MUX al_mux_b0_0_2 (
    .i0(i4),
    .i1(i5),
    .sel(sel[0]),
    .o(B0_2));
  AL_MUX al_mux_b0_0_3 (
    .i0(i6),
    .i1(i7),
    .sel(sel[0]),
    .o(B0_3));
  AL_MUX al_mux_b0_0_4 (
    .i0(i8),
    .i1(i9),
    .sel(sel[0]),
    .o(B0_4));
  AL_MUX al_mux_b0_0_5 (
    .i0(i10),
    .i1(i11),
    .sel(sel[0]),
    .o(B0_5));
  AL_MUX al_mux_b0_0_6 (
    .i0(i12),
    .i1(i13),
    .sel(sel[0]),
    .o(B0_6));
  AL_MUX al_mux_b0_0_7 (
    .i0(i14),
    .i1(i15),
    .sel(sel[0]),
    .o(B0_7));
  AL_MUX al_mux_b0_0_8 (
    .i0(i16),
    .i1(i17),
    .sel(sel[0]),
    .o(B0_8));
  AL_MUX al_mux_b0_0_9 (
    .i0(i18),
    .i1(i19),
    .sel(sel[0]),
    .o(B0_9));
  AL_MUX al_mux_b0_1_0 (
    .i0(B0_0),
    .i1(B0_1),
    .sel(sel[1]),
    .o(B1_0));
  AL_MUX al_mux_b0_1_1 (
    .i0(B0_2),
    .i1(B0_3),
    .sel(sel[1]),
    .o(B1_1));
  AL_MUX al_mux_b0_1_2 (
    .i0(B0_4),
    .i1(B0_5),
    .sel(sel[1]),
    .o(B1_2));
  AL_MUX al_mux_b0_1_3 (
    .i0(B0_6),
    .i1(B0_7),
    .sel(sel[1]),
    .o(B1_3));
  AL_MUX al_mux_b0_1_4 (
    .i0(B0_8),
    .i1(B0_9),
    .sel(sel[1]),
    .o(B1_4));
  AL_MUX al_mux_b0_1_5 (
    .i0(B0_10),
    .i1(B0_11),
    .sel(sel[1]),
    .o(B1_5));
  AL_MUX al_mux_b0_1_6 (
    .i0(B0_12),
    .i1(B0_13),
    .sel(sel[1]),
    .o(B1_6));
  AL_MUX al_mux_b0_1_7 (
    .i0(B0_14),
    .i1(B0_15),
    .sel(sel[1]),
    .o(B1_7));
  AL_MUX al_mux_b0_2_0 (
    .i0(B1_0),
    .i1(B1_1),
    .sel(sel[2]),
    .o(B2_0));
  AL_MUX al_mux_b0_2_1 (
    .i0(B1_2),
    .i1(B1_3),
    .sel(sel[2]),
    .o(B2_1));
  AL_MUX al_mux_b0_2_2 (
    .i0(B1_4),
    .i1(B1_5),
    .sel(sel[2]),
    .o(B2_2));
  AL_MUX al_mux_b0_2_3 (
    .i0(B1_6),
    .i1(B1_7),
    .sel(sel[2]),
    .o(B2_3));
  AL_MUX al_mux_b0_3_0 (
    .i0(B2_0),
    .i1(B2_1),
    .sel(sel[3]),
    .o(B3_0));
  AL_MUX al_mux_b0_3_1 (
    .i0(B2_2),
    .i1(B2_3),
    .sel(sel[3]),
    .o(B3_1));
  AL_MUX al_mux_b0_4_0 (
    .i0(B3_0),
    .i1(B3_1),
    .sel(sel[4]),
    .o(o));

endmodule 

module ne_w1
  (
  i0,
  i1,
  o
  );

  input i0;
  input i1;
  output o;


  xor diff_0 (o, i0, i1);

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

module AL_FADD
  (
  input a,
  input b,
  input c,
  output sum,
  output cout
  );

  wire prop;
  wire not_prop;
  wire sel_i0;
  wire sel_i1;

  xor u0 (prop, a, b);
  xor u1 (sum, prop, c);
  not u2 (not_prop, prop);
  and u3 (sel_i1, prop, c);
  and u4 (sel_i0, not_prop, a);
  or  u5 (cout, sel_i0, sel_i1);

endmodule

